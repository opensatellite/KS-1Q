///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: reboot.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::SmartFusion2> <Die::M2S010> <Package::144 TQ>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module reboot( clk, rst, flag_, port4 );
input port1, port2;
output port3;
inout port4;

//<statements>

endmodule

