`timescale 1 ns/100 ps
// Version: v11.7 11.7.0.119


module MSS_010(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN,
       MMUART0_DCD_MGPIO22B_IN,
       MMUART0_DSR_MGPIO20B_IN,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN,
       MMUART0_RI_MGPIO21B_IN,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN,
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN,
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN,
       SPI1_SCK_IN,
       SPI1_SDI_MGPIO11A_IN,
       SPI1_SDO_MGPIO12A_IN,
       SPI1_SS0_MGPIO13A_IN,
       SPI1_SS1_MGPIO14A_IN,
       SPI1_SS2_MGPIO15A_IN,
       SPI1_SS3_MGPIO16A_IN,
       SPI1_SS4_MGPIO17A_IN,
       SPI1_SS5_MGPIO18A_IN,
       SPI1_SS6_MGPIO23A_IN,
       SPI1_SS7_MGPIO24A_IN,
       USBC_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT,
       MMUART0_DCD_MGPIO22B_OUT,
       MMUART0_DSR_MGPIO20B_OUT,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT,
       MMUART0_RI_MGPIO21B_OUT,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT,
       SPI1_SCK_OUT,
       SPI1_SDI_MGPIO11A_OUT,
       SPI1_SDO_MGPIO12A_OUT,
       SPI1_SS0_MGPIO13A_OUT,
       SPI1_SS1_MGPIO14A_OUT,
       SPI1_SS2_MGPIO15A_OUT,
       SPI1_SS3_MGPIO16A_OUT,
       SPI1_SS4_MGPIO17A_OUT,
       SPI1_SS5_MGPIO18A_OUT,
       SPI1_SS6_MGPIO23A_OUT,
       SPI1_SS7_MGPIO24A_OUT,
       USBC_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE,
       MMUART0_DCD_MGPIO22B_OE,
       MMUART0_DSR_MGPIO20B_OE,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE,
       MMUART0_RI_MGPIO21B_OE,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE,
       SPI1_SCK_OE,
       SPI1_SDI_MGPIO11A_OE,
       SPI1_SDO_MGPIO12A_OE,
       SPI1_SS0_MGPIO13A_OE,
       SPI1_SS1_MGPIO14A_OE,
       SPI1_SS2_MGPIO15A_OE,
       SPI1_SS3_MGPIO16A_OE,
       SPI1_SS4_MGPIO17A_OE,
       SPI1_SS5_MGPIO18A_OE,
       SPI1_SS6_MGPIO23A_OE,
       SPI1_SS7_MGPIO24A_OE,
       USBC_XCLK_OE
    );
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MMUART0_CTS_USBC_DATA7_MGPIO19B_IN;
input  MMUART0_DCD_MGPIO22B_IN;
input  MMUART0_DSR_MGPIO20B_IN;
input  MMUART0_DTR_USBC_DATA6_MGPIO18B_IN;
input  MMUART0_RI_MGPIO21B_IN;
input  MMUART0_RTS_USBC_DATA5_MGPIO17B_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  SPI0_SS1_USBA_DATA5_MGPIO8A_IN;
input  SPI0_SS2_USBA_DATA6_MGPIO9A_IN;
input  SPI0_SS3_USBA_DATA7_MGPIO10A_IN;
input  SPI1_SCK_IN;
input  SPI1_SDI_MGPIO11A_IN;
input  SPI1_SDO_MGPIO12A_IN;
input  SPI1_SS0_MGPIO13A_IN;
input  SPI1_SS1_MGPIO14A_IN;
input  SPI1_SS2_MGPIO15A_IN;
input  SPI1_SS3_MGPIO16A_IN;
input  SPI1_SS4_MGPIO17A_IN;
input  SPI1_SS5_MGPIO18A_IN;
input  SPI1_SS6_MGPIO23A_IN;
input  SPI1_SS7_MGPIO24A_IN;
input  USBC_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT;
output MMUART0_DCD_MGPIO22B_OUT;
output MMUART0_DSR_MGPIO20B_OUT;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT;
output MMUART0_RI_MGPIO21B_OUT;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OUT;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OUT;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OUT;
output SPI1_SCK_OUT;
output SPI1_SDI_MGPIO11A_OUT;
output SPI1_SDO_MGPIO12A_OUT;
output SPI1_SS0_MGPIO13A_OUT;
output SPI1_SS1_MGPIO14A_OUT;
output SPI1_SS2_MGPIO15A_OUT;
output SPI1_SS3_MGPIO16A_OUT;
output SPI1_SS4_MGPIO17A_OUT;
output SPI1_SS5_MGPIO18A_OUT;
output SPI1_SS6_MGPIO23A_OUT;
output SPI1_SS7_MGPIO24A_OUT;
output USBC_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OE;
output MMUART0_DCD_MGPIO22B_OE;
output MMUART0_DSR_MGPIO20B_OE;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OE;
output MMUART0_RI_MGPIO21B_OE;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OE;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OE;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OE;
output SPI1_SCK_OE;
output SPI1_SDI_MGPIO11A_OE;
output SPI1_SDO_MGPIO12A_OE;
output SPI1_SS0_MGPIO13A_OE;
output SPI1_SS1_MGPIO14A_OE;
output SPI1_SS2_MGPIO15A_OE;
output SPI1_SS3_MGPIO16A_OE;
output SPI1_SS4_MGPIO17A_OE;
output SPI1_SS5_MGPIO18A_OE;
output SPI1_SS6_MGPIO23A_OE;
output SPI1_SS7_MGPIO24A_OE;
output USBC_XCLK_OE;

    parameter INIT = 'h0 ;
    parameter ACT_UBITS = 'hFFFFFFFFFFFFFF ;
    parameter MEMORYFILE = "" ;
    parameter RTC_MAIN_XTL_FREQ = 0.0 ;
    parameter RTC_MAIN_XTL_MODE = "1" ;
    parameter DDR_CLK_FREQ = 0.0 ;
    
endmodule


module XTLOSC_FAB(
       A,
       CLKOUT
    );
input  A;
output CLKOUT;

    
endmodule


module XTLOSC(
       XTL,
       CLKOUT
    );
input  XTL;
output CLKOUT;

    parameter MODE = 'h3 ;
    parameter FREQUENCY = 20.0 ;
    
endmodule


module test_4463andcpuopration_MSS(
       CoreAPB3_0_APBmslave3_PADDR,
       CoreAPB3_0_APBmslave3_PWDATA,
       Glue_Logic_0_Flag_Int_0,
       test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       SPI_CLK_c,
       CAN1_RX_c,
       CoreAPB3_0_APBmslave3_PENABLE,
       test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx,
       CoreAPB3_0_APBmslave3_PWRITE,
       SW_c,
       RX_SDN_c,
       Z3V_EN_c,
       L4463_TX_CS_c,
       L4463_RX_CS_c,
       TX_SDN_c,
       L3V3_EN1_c,
       ADC_CSTART_c,
       TXD4_c,
       SPI_FRAM_CS_c,
       SPI_MOSI_c,
       ADC_CS_c,
       ADC_FS_c,
       ADC_PWDN_c,
       L4V_EN_c,
       ANT_SW1_c,
       test_4463andcpuopration_MSS_0_GPIO_15_M2F,
       L3V3_EN2_c,
       CAN1_TX_c,
       N_623_i_0,
       ADC_INT_c,
       L4V_PG_c,
       BOARD_NO_c,
       RXD4_c,
       SPI_MISO_c,
       SYSRESET_0_POWER_ON_RESET_N,
       OSC_0_XTLOSC_O2F
    );
output [31:0] CoreAPB3_0_APBmslave3_PADDR;
output [31:0] CoreAPB3_0_APBmslave3_PWDATA;
input  [0:0] Glue_Logic_0_Flag_Int_0;
input  [31:0] test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA;
output test_4463andcpuopration_MSS_0_GPIO_1_M2F;
output SPI_CLK_c;
output CAN1_RX_c;
output CoreAPB3_0_APBmslave3_PENABLE;
output test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx;
output CoreAPB3_0_APBmslave3_PWRITE;
output SW_c;
output RX_SDN_c;
output Z3V_EN_c;
output L4463_TX_CS_c;
output L4463_RX_CS_c;
output TX_SDN_c;
output L3V3_EN1_c;
output ADC_CSTART_c;
output TXD4_c;
output SPI_FRAM_CS_c;
output SPI_MOSI_c;
output ADC_CS_c;
output ADC_FS_c;
output ADC_PWDN_c;
output L4V_EN_c;
output ANT_SW1_c;
output test_4463andcpuopration_MSS_0_GPIO_15_M2F;
output L3V3_EN2_c;
input  CAN1_TX_c;
input  N_623_i_0;
input  ADC_INT_c;
input  L4V_PG_c;
input  BOARD_NO_c;
input  RXD4_c;
input  SPI_MISO_c;
input  SYSRESET_0_POWER_ON_RESET_N;
input  OSC_0_XTLOSC_O2F;

    wire I2C1_SCL_MGPIO1A_H2F_B, VCC_net_1, GND_net_1;
    
    CLKINT MSS_ADLIB_INST_RNIHTQ8 (.A(I2C1_SCL_MGPIO1A_H2F_B), .Y(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F));
    VCC VCC (.Y(VCC_net_1));
    MSS_010 #( .INIT(1438'h0000000000000030000000000000000000000000000000000000000000000000000000000000000000000000000000000C030000300003000000000000000000000000000000000E00000000F000000000000000000000000000000007FFFFFFFB000001007C33C00000200608D00000003FFFFE00000000000241DC000000F0E01C00000182D754010842108421800001FE34001FF8000000400000000020031007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE(""), .DDR_CLK_FREQ(0.0)
         )  MSS_ADLIB_INST (.CAN_RXBUS_MGPIO3A_H2F_A(), 
        .CAN_RXBUS_MGPIO3A_H2F_B(), .CAN_TX_EBL_MGPIO4A_H2F_A(), 
        .CAN_TX_EBL_MGPIO4A_H2F_B(), .CAN_TXBUS_MGPIO2A_H2F_A(
        CAN1_RX_c), .CAN_TXBUS_MGPIO2A_H2F_B(), .CLK_CONFIG_APB(), 
        .COMMS_INT(), .CONFIG_PRESET_N(), .EDAC_ERROR({nc0, nc1, nc2, 
        nc3, nc4, nc5, nc6, nc7}), .F_FM0_RDATA({nc8, nc9, nc10, nc11, 
        nc12, nc13, nc14, nc15, nc16, nc17, nc18, nc19, nc20, nc21, 
        nc22, nc23, nc24, nc25, nc26, nc27, nc28, nc29, nc30, nc31, 
        nc32, nc33, nc34, nc35, nc36, nc37, nc38, nc39}), 
        .F_FM0_READYOUT(), .F_FM0_RESP(), .F_HM0_ADDR({
        CoreAPB3_0_APBmslave3_PADDR[31], 
        CoreAPB3_0_APBmslave3_PADDR[30], 
        CoreAPB3_0_APBmslave3_PADDR[29], 
        CoreAPB3_0_APBmslave3_PADDR[28], 
        CoreAPB3_0_APBmslave3_PADDR[27], 
        CoreAPB3_0_APBmslave3_PADDR[26], 
        CoreAPB3_0_APBmslave3_PADDR[25], 
        CoreAPB3_0_APBmslave3_PADDR[24], 
        CoreAPB3_0_APBmslave3_PADDR[23], 
        CoreAPB3_0_APBmslave3_PADDR[22], 
        CoreAPB3_0_APBmslave3_PADDR[21], 
        CoreAPB3_0_APBmslave3_PADDR[20], 
        CoreAPB3_0_APBmslave3_PADDR[19], 
        CoreAPB3_0_APBmslave3_PADDR[18], 
        CoreAPB3_0_APBmslave3_PADDR[17], 
        CoreAPB3_0_APBmslave3_PADDR[16], 
        CoreAPB3_0_APBmslave3_PADDR[15], 
        CoreAPB3_0_APBmslave3_PADDR[14], 
        CoreAPB3_0_APBmslave3_PADDR[13], 
        CoreAPB3_0_APBmslave3_PADDR[12], 
        CoreAPB3_0_APBmslave3_PADDR[11], 
        CoreAPB3_0_APBmslave3_PADDR[10], 
        CoreAPB3_0_APBmslave3_PADDR[9], CoreAPB3_0_APBmslave3_PADDR[8], 
        CoreAPB3_0_APBmslave3_PADDR[7], CoreAPB3_0_APBmslave3_PADDR[6], 
        CoreAPB3_0_APBmslave3_PADDR[5], CoreAPB3_0_APBmslave3_PADDR[4], 
        CoreAPB3_0_APBmslave3_PADDR[3], CoreAPB3_0_APBmslave3_PADDR[2], 
        CoreAPB3_0_APBmslave3_PADDR[1], CoreAPB3_0_APBmslave3_PADDR[0]})
        , .F_HM0_ENABLE(CoreAPB3_0_APBmslave3_PENABLE), .F_HM0_SEL(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), 
        .F_HM0_SIZE({nc40, nc41}), .F_HM0_TRANS1(), .F_HM0_WDATA({
        CoreAPB3_0_APBmslave3_PWDATA[31], 
        CoreAPB3_0_APBmslave3_PWDATA[30], 
        CoreAPB3_0_APBmslave3_PWDATA[29], 
        CoreAPB3_0_APBmslave3_PWDATA[28], 
        CoreAPB3_0_APBmslave3_PWDATA[27], 
        CoreAPB3_0_APBmslave3_PWDATA[26], 
        CoreAPB3_0_APBmslave3_PWDATA[25], 
        CoreAPB3_0_APBmslave3_PWDATA[24], 
        CoreAPB3_0_APBmslave3_PWDATA[23], 
        CoreAPB3_0_APBmslave3_PWDATA[22], 
        CoreAPB3_0_APBmslave3_PWDATA[21], 
        CoreAPB3_0_APBmslave3_PWDATA[20], 
        CoreAPB3_0_APBmslave3_PWDATA[19], 
        CoreAPB3_0_APBmslave3_PWDATA[18], 
        CoreAPB3_0_APBmslave3_PWDATA[17], 
        CoreAPB3_0_APBmslave3_PWDATA[16], 
        CoreAPB3_0_APBmslave3_PWDATA[15], 
        CoreAPB3_0_APBmslave3_PWDATA[14], 
        CoreAPB3_0_APBmslave3_PWDATA[13], 
        CoreAPB3_0_APBmslave3_PWDATA[12], 
        CoreAPB3_0_APBmslave3_PWDATA[11], 
        CoreAPB3_0_APBmslave3_PWDATA[10], 
        CoreAPB3_0_APBmslave3_PWDATA[9], 
        CoreAPB3_0_APBmslave3_PWDATA[8], 
        CoreAPB3_0_APBmslave3_PWDATA[7], 
        CoreAPB3_0_APBmslave3_PWDATA[6], 
        CoreAPB3_0_APBmslave3_PWDATA[5], 
        CoreAPB3_0_APBmslave3_PWDATA[4], 
        CoreAPB3_0_APBmslave3_PWDATA[3], 
        CoreAPB3_0_APBmslave3_PWDATA[2], 
        CoreAPB3_0_APBmslave3_PWDATA[1], 
        CoreAPB3_0_APBmslave3_PWDATA[0]}), .F_HM0_WRITE(
        CoreAPB3_0_APBmslave3_PWRITE), .FAB_CHRGVBUS(), 
        .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), .FAB_DPPULLDOWN(), 
        .FAB_DRVVBUS(), .FAB_IDPULLUP(), .FAB_OPMODE({nc42, nc43}), 
        .FAB_SUSPENDM(), .FAB_TERMSEL(), .FAB_TXVALID(), .FAB_VCONTROL({
        nc44, nc45, nc46, nc47}), .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({
        nc48, nc49}), .FAB_XDATAOUT({nc50, nc51, nc52, nc53, nc54, 
        nc55, nc56, nc57}), .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc58, 
        nc59}), .FIC32_1_MASTER({nc60, nc61}), .FPGA_RESET_N(), 
        .GTX_CLK(), .H2F_INTERRUPT({nc62, nc63, nc64, nc65, nc66, nc67, 
        nc68, nc69, nc70, nc71, nc72, nc73, nc74, nc75, nc76, nc77}), 
        .H2F_NMI(), .H2FCALIB(), .I2C0_SCL_MGPIO31B_H2F_A(), 
        .I2C0_SCL_MGPIO31B_H2F_B(), .I2C0_SDA_MGPIO30B_H2F_A(), 
        .I2C0_SDA_MGPIO30B_H2F_B(), .I2C1_SCL_MGPIO1A_H2F_A(), 
        .I2C1_SCL_MGPIO1A_H2F_B(I2C1_SCL_MGPIO1A_H2F_B), 
        .I2C1_SDA_MGPIO0A_H2F_A(), .I2C1_SDA_MGPIO0A_H2F_B(SW_c), 
        .MDCF(), .MDOENF(), .MDOF(), .MMUART0_CTS_MGPIO19B_H2F_A(), 
        .MMUART0_CTS_MGPIO19B_H2F_B(RX_SDN_c), 
        .MMUART0_DCD_MGPIO22B_H2F_A(), .MMUART0_DCD_MGPIO22B_H2F_B(
        Z3V_EN_c), .MMUART0_DSR_MGPIO20B_H2F_A(), 
        .MMUART0_DSR_MGPIO20B_H2F_B(L4463_TX_CS_c), 
        .MMUART0_DTR_MGPIO18B_H2F_A(), .MMUART0_DTR_MGPIO18B_H2F_B(
        L4463_RX_CS_c), .MMUART0_RI_MGPIO21B_H2F_A(), 
        .MMUART0_RI_MGPIO21B_H2F_B(TX_SDN_c), 
        .MMUART0_RTS_MGPIO17B_H2F_A(), .MMUART0_RTS_MGPIO17B_H2F_B(
        L3V3_EN1_c), .MMUART0_RXD_MGPIO28B_H2F_A(), 
        .MMUART0_RXD_MGPIO28B_H2F_B(), .MMUART0_SCK_MGPIO29B_H2F_A(), 
        .MMUART0_SCK_MGPIO29B_H2F_B(ADC_CSTART_c), 
        .MMUART0_TXD_MGPIO27B_H2F_A(TXD4_c), 
        .MMUART0_TXD_MGPIO27B_H2F_B(), .MMUART1_DTR_MGPIO12B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_B(), 
        .MMUART1_RXD_MGPIO26B_H2F_A(), .MMUART1_RXD_MGPIO26B_H2F_B(), 
        .MMUART1_SCK_MGPIO25B_H2F_A(), .MMUART1_SCK_MGPIO25B_H2F_B(
        SPI_FRAM_CS_c), .MMUART1_TXD_MGPIO24B_H2F_A(), 
        .MMUART1_TXD_MGPIO24B_H2F_B(), .MPLL_LOCK(), 
        .PER2_FABRIC_PADDR({nc78, nc79, nc80, nc81, nc82, nc83, nc84, 
        nc85, nc86, nc87, nc88, nc89, nc90, nc91}), 
        .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc92, nc93, nc94, nc95, nc96, nc97, nc98, 
        nc99, nc100, nc101, nc102, nc103, nc104, nc105, nc106, nc107, 
        nc108, nc109, nc110, nc111, nc112, nc113, nc114, nc115, nc116, 
        nc117, nc118, nc119, nc120, nc121, nc122, nc123}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(SPI_CLK_c), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(SPI_MOSI_c), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(ADC_CS_c), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(ADC_FS_c), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(
        ADC_PWDN_c), .SPI0_SS4_MGPIO19A_H2F_A(), 
        .SPI0_SS5_MGPIO20A_H2F_A(), .SPI0_SS6_MGPIO21A_H2F_A(), 
        .SPI0_SS7_MGPIO22A_H2F_A(), .SPI1_CLK_OUT(), 
        .SPI1_SDI_MGPIO11A_H2F_A(), .SPI1_SDI_MGPIO11A_H2F_B(), 
        .SPI1_SDO_MGPIO12A_H2F_A(), .SPI1_SDO_MGPIO12A_H2F_B(L4V_EN_c), 
        .SPI1_SS0_MGPIO13A_H2F_A(), .SPI1_SS0_MGPIO13A_H2F_B(ANT_SW1_c)
        , .SPI1_SS1_MGPIO14A_H2F_A(), .SPI1_SS1_MGPIO14A_H2F_B(), 
        .SPI1_SS2_MGPIO15A_H2F_A(), .SPI1_SS2_MGPIO15A_H2F_B(
        test_4463andcpuopration_MSS_0_GPIO_15_M2F), 
        .SPI1_SS3_MGPIO16A_H2F_A(), .SPI1_SS3_MGPIO16A_H2F_B(
        L3V3_EN2_c), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc124, nc125, nc126, nc127, 
        nc128, nc129, nc130, nc131, nc132, nc133}), .TRACECLK(), 
        .TRACEDATA({nc134, nc135, nc136, nc137}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc138, nc139, nc140, 
        nc141}), .TXDF({nc142, nc143, nc144, nc145, nc146, nc147, 
        nc148, nc149}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc150, nc151, nc152, nc153})
        , .F_BRESP_HRESP0({nc154, nc155}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc156, nc157, nc158, nc159, nc160, nc161, 
        nc162, nc163, nc164, nc165, nc166, nc167, nc168, nc169, nc170, 
        nc171, nc172, nc173, nc174, nc175, nc176, nc177, nc178, nc179, 
        nc180, nc181, nc182, nc183, nc184, nc185, nc186, nc187, nc188, 
        nc189, nc190, nc191, nc192, nc193, nc194, nc195, nc196, nc197, 
        nc198, nc199, nc200, nc201, nc202, nc203, nc204, nc205, nc206, 
        nc207, nc208, nc209, nc210, nc211, nc212, nc213, nc214, nc215, 
        nc216, nc217, nc218, nc219}), .F_RID({nc220, nc221, nc222, 
        nc223}), .F_RLAST(), .F_RRESP_HRESP1({nc224, nc225}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc226, nc227, 
        nc228, nc229, nc230, nc231, nc232, nc233, nc234, nc235, nc236, 
        nc237, nc238, nc239, nc240, nc241}), .MDDR_FABRIC_PREADY(), 
        .MDDR_FABRIC_PSLVERR(), .CAN_RXBUS_F2H_SCP(CAN1_TX_c), 
        .CAN_TX_EBL_F2H_SCP(VCC_net_1), .CAN_TXBUS_F2H_SCP(VCC_net_1), 
        .COLF(VCC_net_1), .CRSF(VCC_net_1), .F2_DMAREADY({VCC_net_1, 
        VCC_net_1}), .F2H_INTERRUPT({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, Glue_Logic_0_Flag_Int_0[0]}), .F2HCALIB(
        VCC_net_1), .F_DMAREADY({VCC_net_1, VCC_net_1}), .F_FM0_ADDR({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_FM0_ENABLE(GND_net_1), 
        .F_FM0_MASTLOCK(GND_net_1), .F_FM0_READY(VCC_net_1), 
        .F_FM0_SEL(GND_net_1), .F_FM0_SIZE({GND_net_1, GND_net_1}), 
        .F_FM0_TRANS1(GND_net_1), .F_FM0_WDATA({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_FM0_WRITE(GND_net_1), .F_HM0_RDATA({
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[31], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[30], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[29], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[28], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[27], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[26], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[25], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[24], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[23], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[22], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[21], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[20], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[19], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[18], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[17], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[16], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[15], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[14], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[13], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[12], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[11], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[10], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[9], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[8], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[7], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[6], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[5], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[4], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[3], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[2], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[1], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[0]}), 
        .F_HM0_READY(N_623_i_0), .F_HM0_RESP(GND_net_1), .FAB_AVALID(
        VCC_net_1), .FAB_HOSTDISCON(VCC_net_1), .FAB_IDDIG(VCC_net_1), 
        .FAB_LINESTATE({VCC_net_1, VCC_net_1}), .FAB_M3_RESET_N(
        VCC_net_1), .FAB_PLL_LOCK(VCC_net_1), .FAB_RXACTIVE(VCC_net_1), 
        .FAB_RXERROR(VCC_net_1), .FAB_RXVALID(VCC_net_1), 
        .FAB_RXVALIDH(GND_net_1), .FAB_SESSEND(VCC_net_1), 
        .FAB_TXREADY(VCC_net_1), .FAB_VBUSVALID(VCC_net_1), 
        .FAB_VSTATUS({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), .FAB_XDATAIN({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .GTX_CLKPF(VCC_net_1), 
        .I2C0_BCLK(VCC_net_1), .I2C0_SCL_F2H_SCP(VCC_net_1), 
        .I2C0_SDA_F2H_SCP(VCC_net_1), .I2C1_BCLK(VCC_net_1), 
        .I2C1_SCL_F2H_SCP(VCC_net_1), .I2C1_SDA_F2H_SCP(VCC_net_1), 
        .MDIF(VCC_net_1), .MGPIO0A_F2H_GPIN(VCC_net_1), 
        .MGPIO10A_F2H_GPIN(VCC_net_1), .MGPIO11A_F2H_GPIN(VCC_net_1), 
        .MGPIO11B_F2H_GPIN(VCC_net_1), .MGPIO12A_F2H_GPIN(VCC_net_1), 
        .MGPIO13A_F2H_GPIN(VCC_net_1), .MGPIO14A_F2H_GPIN(VCC_net_1), 
        .MGPIO15A_F2H_GPIN(VCC_net_1), .MGPIO16A_F2H_GPIN(VCC_net_1), 
        .MGPIO17B_F2H_GPIN(VCC_net_1), .MGPIO18B_F2H_GPIN(VCC_net_1), 
        .MGPIO19B_F2H_GPIN(VCC_net_1), .MGPIO1A_F2H_GPIN(VCC_net_1), 
        .MGPIO20B_F2H_GPIN(VCC_net_1), .MGPIO21B_F2H_GPIN(VCC_net_1), 
        .MGPIO22B_F2H_GPIN(VCC_net_1), .MGPIO24B_F2H_GPIN(VCC_net_1), 
        .MGPIO25B_F2H_GPIN(VCC_net_1), .MGPIO26B_F2H_GPIN(ADC_INT_c), 
        .MGPIO27B_F2H_GPIN(GND_net_1), .MGPIO28B_F2H_GPIN(GND_net_1), 
        .MGPIO29B_F2H_GPIN(VCC_net_1), .MGPIO2A_F2H_GPIN(VCC_net_1), 
        .MGPIO30B_F2H_GPIN(L4V_PG_c), .MGPIO31B_F2H_GPIN(BOARD_NO_c), 
        .MGPIO3A_F2H_GPIN(VCC_net_1), .MGPIO4A_F2H_GPIN(VCC_net_1), 
        .MGPIO5A_F2H_GPIN(VCC_net_1), .MGPIO6A_F2H_GPIN(VCC_net_1), 
        .MGPIO7A_F2H_GPIN(VCC_net_1), .MGPIO8A_F2H_GPIN(VCC_net_1), 
        .MGPIO9A_F2H_GPIN(VCC_net_1), .MMUART0_CTS_F2H_SCP(VCC_net_1), 
        .MMUART0_DCD_F2H_SCP(VCC_net_1), .MMUART0_DSR_F2H_SCP(
        VCC_net_1), .MMUART0_DTR_F2H_SCP(VCC_net_1), 
        .MMUART0_RI_F2H_SCP(VCC_net_1), .MMUART0_RTS_F2H_SCP(VCC_net_1)
        , .MMUART0_RXD_F2H_SCP(RXD4_c), .MMUART0_SCK_F2H_SCP(VCC_net_1)
        , .MMUART0_TXD_F2H_SCP(VCC_net_1), .MMUART1_CTS_F2H_SCP(
        VCC_net_1), .MMUART1_DCD_F2H_SCP(VCC_net_1), 
        .MMUART1_DSR_F2H_SCP(VCC_net_1), .MMUART1_RI_F2H_SCP(VCC_net_1)
        , .MMUART1_RTS_F2H_SCP(VCC_net_1), .MMUART1_RXD_F2H_SCP(
        VCC_net_1), .MMUART1_SCK_F2H_SCP(VCC_net_1), 
        .MMUART1_TXD_F2H_SCP(VCC_net_1), .PER2_FABRIC_PRDATA({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1}), .PER2_FABRIC_PREADY(VCC_net_1), 
        .PER2_FABRIC_PSLVERR(VCC_net_1), .RCGF({VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .RX_CLKPF(VCC_net_1), 
        .RX_DVF(VCC_net_1), .RX_ERRF(VCC_net_1), .RX_EV(VCC_net_1), 
        .RXDF({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .SLEEPHOLDREQ(GND_net_1), 
        .SMBALERT_NI0(VCC_net_1), .SMBALERT_NI1(VCC_net_1), 
        .SMBSUS_NI0(VCC_net_1), .SMBSUS_NI1(VCC_net_1), .SPI0_CLK_IN(
        SPI_CLK_c), .SPI0_SDI_F2H_SCP(SPI_MISO_c), .SPI0_SDO_F2H_SCP(
        VCC_net_1), .SPI0_SS0_F2H_SCP(VCC_net_1), .SPI0_SS1_F2H_SCP(
        VCC_net_1), .SPI0_SS2_F2H_SCP(VCC_net_1), .SPI0_SS3_F2H_SCP(
        VCC_net_1), .SPI1_CLK_IN(VCC_net_1), .SPI1_SDI_F2H_SCP(
        VCC_net_1), .SPI1_SDO_F2H_SCP(VCC_net_1), .SPI1_SS0_F2H_SCP(
        VCC_net_1), .SPI1_SS1_F2H_SCP(VCC_net_1), .SPI1_SS2_F2H_SCP(
        VCC_net_1), .SPI1_SS3_F2H_SCP(VCC_net_1), .TX_CLKPF(VCC_net_1), 
        .USER_MSS_GPIO_RESET_N(VCC_net_1), .USER_MSS_RESET_N(
        SYSRESET_0_POWER_ON_RESET_N), .XCLK_FAB(VCC_net_1), .CLK_BASE(
        OSC_0_XTLOSC_O2F), .CLK_MDDR_APB(VCC_net_1), .F_ARADDR_HADDR1({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1}), .F_ARBURST_HTRANS1({GND_net_1, 
        GND_net_1}), .F_ARID_HSEL1({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_ARLEN_HBURST1({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_ARLOCK_HMASTLOCK1({GND_net_1, GND_net_1}), 
        .F_ARSIZE_HSIZE1({GND_net_1, GND_net_1}), .F_ARVALID_HWRITE1(
        GND_net_1), .F_AWADDR_HADDR0({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .F_AWBURST_HTRANS0({GND_net_1, GND_net_1}), .F_AWID_HSEL0({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .F_AWLEN_HBURST0({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLOCK_HMASTLOCK0({GND_net_1, GND_net_1}), .F_AWSIZE_HSIZE0({
        GND_net_1, GND_net_1}), .F_AWVALID_HWRITE0(GND_net_1), 
        .F_BREADY(GND_net_1), .F_RMW_AXI(GND_net_1), .F_RREADY(
        GND_net_1), .F_WDATA_HWDATA01({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_WID_HREADY01({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_WLAST(GND_net_1), .F_WSTRB({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_WVALID(GND_net_1), 
        .FPGA_MDDR_ARESET_N(VCC_net_1), .MDDR_FABRIC_PADDR({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .MDDR_FABRIC_PENABLE(
        VCC_net_1), .MDDR_FABRIC_PSEL(VCC_net_1), .MDDR_FABRIC_PWDATA({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .MDDR_FABRIC_PWRITE(VCC_net_1), .PRESET_N(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND_net_1), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND_net_1), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND_net_1), .DM_IN({GND_net_1, 
        GND_net_1, GND_net_1}), .DRAM_DQ_IN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .DRAM_DQS_IN({GND_net_1, GND_net_1, GND_net_1}), 
        .DRAM_FIFO_WE_IN({GND_net_1, GND_net_1}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND_net_1), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND_net_1), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND_net_1), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND_net_1), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND_net_1), 
        .MMUART0_DCD_MGPIO22B_IN(GND_net_1), .MMUART0_DSR_MGPIO20B_IN(
        GND_net_1), .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND_net_1), 
        .MMUART0_RI_MGPIO21B_IN(GND_net_1), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND_net_1), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(GND_net_1), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND_net_1), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND_net_1), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(GND_net_1), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND_net_1), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND_net_1), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND_net_1), 
        .RGMII_MDC_RMII_MDC_IN(GND_net_1), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND_net_1), 
        .RGMII_RX_CLK_IN(GND_net_1), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND_net_1), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND_net_1), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND_net_1), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND_net_1), 
        .RGMII_RXD3_USBB_DATA4_IN(GND_net_1), .RGMII_TX_CLK_IN(
        GND_net_1), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND_net_1), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND_net_1), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND_net_1), 
        .RGMII_TXD2_USBB_DATA5_IN(GND_net_1), 
        .RGMII_TXD3_USBB_DATA6_IN(GND_net_1), .SPI0_SCK_USBA_XCLK_IN(
        GND_net_1), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(GND_net_1), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND_net_1), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(GND_net_1), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND_net_1), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND_net_1), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND_net_1), .SPI1_SCK_IN(
        GND_net_1), .SPI1_SDI_MGPIO11A_IN(GND_net_1), 
        .SPI1_SDO_MGPIO12A_IN(GND_net_1), .SPI1_SS0_MGPIO13A_IN(
        GND_net_1), .SPI1_SS1_MGPIO14A_IN(GND_net_1), 
        .SPI1_SS2_MGPIO15A_IN(GND_net_1), .SPI1_SS3_MGPIO16A_IN(
        GND_net_1), .SPI1_SS4_MGPIO17A_IN(GND_net_1), 
        .SPI1_SS5_MGPIO18A_IN(GND_net_1), .SPI1_SS6_MGPIO23A_IN(
        GND_net_1), .SPI1_SS7_MGPIO24A_IN(GND_net_1), .USBC_XCLK_IN(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({nc242, nc243, 
        nc244, nc245, nc246, nc247, nc248, nc249, nc250, nc251, nc252, 
        nc253, nc254, nc255, nc256, nc257}), .DRAM_BA({nc258, nc259, 
        nc260}), .DRAM_CASN(), .DRAM_CKE(), .DRAM_CLK(), .DRAM_CSN(), 
        .DRAM_DM_RDQS_OUT({nc261, nc262, nc263}), .DRAM_DQ_OUT({nc264, 
        nc265, nc266, nc267, nc268, nc269, nc270, nc271, nc272, nc273, 
        nc274, nc275, nc276, nc277, nc278, nc279, nc280, nc281}), 
        .DRAM_DQS_OUT({nc282, nc283, nc284}), .DRAM_FIFO_WE_OUT({nc285, 
        nc286}), .DRAM_ODT(), .DRAM_RASN(), .DRAM_RSTN(), .DRAM_WEN(), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(), .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI1_SCK_OUT(), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(), 
        .SPI1_SS0_MGPIO13A_OUT(), .SPI1_SS1_MGPIO14A_OUT(), 
        .SPI1_SS2_MGPIO15A_OUT(), .SPI1_SS3_MGPIO16A_OUT(), 
        .SPI1_SS4_MGPIO17A_OUT(), .SPI1_SS5_MGPIO18A_OUT(), 
        .SPI1_SS6_MGPIO23A_OUT(), .SPI1_SS7_MGPIO24A_OUT(), 
        .USBC_XCLK_OUT(), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc287, nc288, 
        nc289}), .DRAM_DQ_OE({nc290, nc291, nc292, nc293, nc294, nc295, 
        nc296, nc297, nc298, nc299, nc300, nc301, nc302, nc303, nc304, 
        nc305, nc306, nc307}), .DRAM_DQS_OE({nc308, nc309, nc310}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        ), .SPI0_SS0_USBA_NXT_MGPIO7A_OE(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI1_SCK_OE(), 
        .SPI1_SDI_MGPIO11A_OE(), .SPI1_SDO_MGPIO12A_OE(), 
        .SPI1_SS0_MGPIO13A_OE(), .SPI1_SS1_MGPIO14A_OE(), 
        .SPI1_SS2_MGPIO15A_OE(), .SPI1_SS3_MGPIO16A_OE(), 
        .SPI1_SS4_MGPIO17A_OE(), .SPI1_SS5_MGPIO18A_OE(), 
        .SPI1_SS6_MGPIO23A_OE(), .SPI1_SS7_MGPIO24A_OE(), 
        .USBC_XCLK_OE());
    GND GND (.Y(GND_net_1));
    
endmodule


module Switch(
       stream,
       pn_reg,
       Switch_0_EnOut,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       P_CLK,
       c_in,
       ASM_OUT,
       S_OUT_0,
       P_OUT
    );
input  [0:0] stream;
input  [0:0] pn_reg;
output Switch_0_EnOut;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  P_CLK;
output c_in;
input  ASM_OUT;
input  S_OUT_0;
input  P_OUT;

    wire VCC_net_1, EnOut_2_net_1, GND_net_1, Out_4, N_118;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'hB) )  EnOut_2 (.A(S_OUT_0), .B(stream[0]), .Y(
        EnOut_2_net_1));
    SLE EnOut (.D(EnOut_2_net_1), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Switch_0_EnOut));
    CFG4 #( .INIT(16'h4EE4) )  Out_4_u (.A(S_OUT_0), .B(N_118), .C(
        P_OUT), .D(pn_reg[0]), .Y(Out_4));
    CFG2 #( .INIT(4'h4) )  Out_4_0 (.A(stream[0]), .B(ASM_OUT), .Y(
        N_118));
    SLE Out (.D(Out_4), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(c_in));
    
endmodule


module CPU_W_HDL_R(
       CPU_W_HDL_R_0_TM_Packet_Counter,
       CPU_W_HDL_R_0_USER_RA_TRP1_9,
       CPU_W_HDL_R_0_USER_RA_TRP1_0,
       CPU_W_HDL_R_0_USER_RA_TRP1_1,
       CPU_W_HDL_R_0_USER_RA_TRP1_2,
       CPU_W_HDL_R_0_USER_RA_TRP1_3,
       CPU_W_HDL_R_0_USER_RA_TRP1_4,
       CPU_W_HDL_R_0_USER_RA_TRP1_5,
       CPU_W_HDL_R_0_USER_RA_TRP1_6,
       CPU_W_HDL_R_0_USER_RA_TRP1_7,
       ENASM,
       ENASM_i_0,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       P_CLK,
       CPU_W_HDL_R_0_USER_REN_TRP1,
       CPU_W_HDL_R_0_Flag_B_Tx_Finish,
       CPU_W_HDL_R_0_Flag_A_Tx_Finish,
       ENCRC,
       Glue_Logic_0_Flag_B_Tx,
       TXD4_net_0,
       pending,
       En_read_buff
    );
output [31:0] CPU_W_HDL_R_0_TM_Packet_Counter;
output CPU_W_HDL_R_0_USER_RA_TRP1_9;
output CPU_W_HDL_R_0_USER_RA_TRP1_0;
output CPU_W_HDL_R_0_USER_RA_TRP1_1;
output CPU_W_HDL_R_0_USER_RA_TRP1_2;
output CPU_W_HDL_R_0_USER_RA_TRP1_3;
output CPU_W_HDL_R_0_USER_RA_TRP1_4;
output CPU_W_HDL_R_0_USER_RA_TRP1_5;
output CPU_W_HDL_R_0_USER_RA_TRP1_6;
output CPU_W_HDL_R_0_USER_RA_TRP1_7;
output ENASM;
output ENASM_i_0;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  P_CLK;
output CPU_W_HDL_R_0_USER_REN_TRP1;
output CPU_W_HDL_R_0_Flag_B_Tx_Finish;
output CPU_W_HDL_R_0_Flag_A_Tx_Finish;
output ENCRC;
input  Glue_Logic_0_Flag_B_Tx;
input  TXD4_net_0;
input  pending;
input  En_read_buff;

    wire \clock_dec[0]_net_1 , \clock_dec_i_0[0] , 
        \ASM_Count[2]_net_1 , VCC_net_1, N_459_i_0, GND_net_1, 
        \ASM_Count[3]_net_1 , N_458_i_0, \clock_dec[1]_net_1 , 
        \clock_dec_RNO[1]_net_1 , \clock_dec[2]_net_1 , N_103_i_i_0, 
        \Flag_Type[0]_net_1 , Flag_Type11, un1_Flag_B_Tx_Finish17_i_0, 
        \Flag_Type[1]_net_1 , Flag_Type11_i_0, \ASM_Count[0]_net_1 , 
        N_461_i_0, \ASM_Count[1]_net_1 , N_460_i_0, \State[1]_net_1 , 
        \State_ns[1] , N_1296_i_0, Addr, N_136_i_0, N_456_i_0, 
        N_31_i_0, N_3_i_0, Flag_B_Tx_Finish_3, Flag_A_Tx_Finish_3, 
        N_457_i_0, N_29_i_1, pos1_En_ASG_net_1, \Addr_s[0] , N_5_i_0, 
        \Addr_s[1] , \Addr_s[2] , \Addr_s[3] , \Addr_s[4] , 
        \Addr_s[5] , \Addr_s[6] , \Addr_s[7]_net_1 , 
        \TM_Packet_Counter_s[0] , \TM_Packet_Counter_s[1] , 
        \TM_Packet_Counter_s[2] , \TM_Packet_Counter_s[3] , 
        \TM_Packet_Counter_s[4] , \TM_Packet_Counter_s[5] , 
        \TM_Packet_Counter_s[6] , \TM_Packet_Counter_s[7] , 
        \TM_Packet_Counter_s[8] , \TM_Packet_Counter_s[9] , 
        \TM_Packet_Counter_s[10] , \TM_Packet_Counter_s[11] , 
        \TM_Packet_Counter_s[12] , \TM_Packet_Counter_s[13] , 
        \TM_Packet_Counter_s[14] , \TM_Packet_Counter_s[15] , 
        \TM_Packet_Counter_s[16] , \TM_Packet_Counter_s[17] , 
        \TM_Packet_Counter_s[18] , \TM_Packet_Counter_s[19] , 
        \TM_Packet_Counter_s[20] , \TM_Packet_Counter_s[21] , 
        \TM_Packet_Counter_s[22] , \TM_Packet_Counter_s[23] , 
        \TM_Packet_Counter_s[24] , \TM_Packet_Counter_s[25] , 
        \TM_Packet_Counter_s[26] , \TM_Packet_Counter_s[27] , 
        \TM_Packet_Counter_s[28] , \TM_Packet_Counter_s[29] , 
        \TM_Packet_Counter_s[30] , \TM_Packet_Counter_s[31]_net_1 , 
        TM_Packet_Counter_cry_cy, \TM_Packet_Counter_cry[0]_net_1 , 
        \TM_Packet_Counter_cry[1]_net_1 , 
        \TM_Packet_Counter_cry[2]_net_1 , 
        \TM_Packet_Counter_cry[3]_net_1 , 
        \TM_Packet_Counter_cry[4]_net_1 , 
        \TM_Packet_Counter_cry[5]_net_1 , 
        \TM_Packet_Counter_cry[6]_net_1 , 
        \TM_Packet_Counter_cry[7]_net_1 , 
        \TM_Packet_Counter_cry[8]_net_1 , 
        \TM_Packet_Counter_cry[9]_net_1 , 
        \TM_Packet_Counter_cry[10]_net_1 , 
        \TM_Packet_Counter_cry[11]_net_1 , 
        \TM_Packet_Counter_cry[12]_net_1 , 
        \TM_Packet_Counter_cry[13]_net_1 , 
        \TM_Packet_Counter_cry[14]_net_1 , 
        \TM_Packet_Counter_cry[15]_net_1 , 
        \TM_Packet_Counter_cry[16]_net_1 , 
        \TM_Packet_Counter_cry[17]_net_1 , 
        \TM_Packet_Counter_cry[18]_net_1 , 
        \TM_Packet_Counter_cry[19]_net_1 , 
        \TM_Packet_Counter_cry[20]_net_1 , 
        \TM_Packet_Counter_cry[21]_net_1 , 
        \TM_Packet_Counter_cry[22]_net_1 , 
        \TM_Packet_Counter_cry[23]_net_1 , 
        \TM_Packet_Counter_cry[24]_net_1 , 
        \TM_Packet_Counter_cry[25]_net_1 , 
        \TM_Packet_Counter_cry[26]_net_1 , 
        \TM_Packet_Counter_cry[27]_net_1 , 
        \TM_Packet_Counter_cry[28]_net_1 , 
        \TM_Packet_Counter_cry[29]_net_1 , 
        \TM_Packet_Counter_cry[30]_net_1 , Addr_s_366_FCO, 
        \Addr_cry[0]_net_1 , \Addr_cry[1]_net_1 , \Addr_cry[2]_net_1 , 
        \Addr_cry[3]_net_1 , \Addr_cry[4]_net_1 , \Addr_cry[5]_net_1 , 
        \Addr_cry[6]_net_1 , N_1300, N_1292, 
        Flag_B_Tx_Finish_3_f0_0_0_a2_0_0_net_1, N_1288, N_85, N_1366, 
        N_1346_4, N_1287, N_1340, N_1310, N_1343, 
        un1_Flag_B_Tx_Finish17_2_i_i_0_1;
    
    CFG3 #( .INIT(8'h73) )  \Flag_Type_RNO[1]  (.A(N_1292), .B(
        TXD4_net_0), .C(Glue_Logic_0_Flag_B_Tx), .Y(Flag_Type11_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[24]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[24]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[23]_net_1 ), .S(
        \TM_Packet_Counter_s[24] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[24]_net_1 ));
    SLE pos1_En_ASG (.D(ENASM), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pos1_En_ASG_net_1));
    ARI1 #( .INIT(20'h48800) )  \Addr_cry[0]  (.A(VCC_net_1), .B(Addr), 
        .C(CPU_W_HDL_R_0_USER_RA_TRP1_0), .D(GND_net_1), .FCI(
        Addr_s_366_FCO), .S(\Addr_s[0] ), .Y(), .FCO(
        \Addr_cry[0]_net_1 ));
    SLE Flag_A_Tx_Finish (.D(Flag_A_Tx_Finish_3), .CLK(P_CLK), .EN(
        N_1296_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CPU_W_HDL_R_0_Flag_A_Tx_Finish));
    SLE \Addr[6]  (.D(\Addr_s[6] ), .CLK(P_CLK), .EN(N_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_USER_RA_TRP1_6));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[19]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[19]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[18]_net_1 ), .S(
        \TM_Packet_Counter_s[19] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[19]_net_1 ));
    SLE \TM_Packet_Counter[0]  (.D(\TM_Packet_Counter_s[0] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[0]));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[26]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[26]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[25]_net_1 ), .S(
        \TM_Packet_Counter_s[26] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[26]_net_1 ));
    SLE \TM_Packet_Counter[1]  (.D(\TM_Packet_Counter_s[1] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[1]));
    CFG4 #( .INIT(16'hCE00) )  \ASM_Count_RNO[3]  (.A(
        \ASM_Count[2]_net_1 ), .B(\ASM_Count[3]_net_1 ), .C(N_85), .D(
        ENCRC), .Y(N_458_i_0));
    CFG4 #( .INIT(16'hCC4C) )  \Flag_Type_RNI6EBH[0]  (.A(
        Glue_Logic_0_Flag_B_Tx), .B(TXD4_net_0), .C(
        \Flag_Type[0]_net_1 ), .D(\Flag_Type[1]_net_1 ), .Y(
        Flag_Type11));
    ARI1 #( .INIT(20'h48800) )  \Addr_cry[1]  (.A(VCC_net_1), .B(Addr), 
        .C(CPU_W_HDL_R_0_USER_RA_TRP1_1), .D(GND_net_1), .FCI(
        \Addr_cry[0]_net_1 ), .S(\Addr_s[1] ), .Y(), .FCO(
        \Addr_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \Addr_cry[3]  (.A(VCC_net_1), .B(Addr), 
        .C(CPU_W_HDL_R_0_USER_RA_TRP1_3), .D(GND_net_1), .FCI(
        \Addr_cry[2]_net_1 ), .S(\Addr_s[3] ), .Y(), .FCO(
        \Addr_cry[3]_net_1 ));
    CFG4 #( .INIT(16'hF9F0) )  \State_ns_0_0[1]  (.A(
        \Flag_Type[0]_net_1 ), .B(\Flag_Type[1]_net_1 ), .C(N_1340), 
        .D(\State[1]_net_1 ), .Y(\State_ns[1] ));
    SLE \TM_Packet_Counter[29]  (.D(\TM_Packet_Counter_s[29] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[29]));
    ARI1 #( .INIT(20'h48800) )  \Addr_cry[6]  (.A(VCC_net_1), .B(Addr), 
        .C(CPU_W_HDL_R_0_USER_RA_TRP1_6), .D(GND_net_1), .FCI(
        \Addr_cry[5]_net_1 ), .S(\Addr_s[6] ), .Y(), .FCO(
        \Addr_cry[6]_net_1 ));
    CFG4 #( .INIT(16'h020A) )  En_ASG_RNO (.A(ENCRC), .B(
        \State[1]_net_1 ), .C(N_1300), .D(N_1296_i_0), .Y(N_29_i_1));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[8]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[8]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[7]_net_1 ), .S(\TM_Packet_Counter_s[8] )
        , .Y(), .FCO(\TM_Packet_Counter_cry[8]_net_1 ));
    SLE \TM_Packet_Counter[2]  (.D(\TM_Packet_Counter_s[2] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[2]));
    CFG2 #( .INIT(4'h4) )  Flag_B_Tx_Finish_3_f0_0_0_a2_0_0 (.A(
        \Flag_Type[0]_net_1 ), .B(\Flag_Type[1]_net_1 ), .Y(
        Flag_B_Tx_Finish_3_f0_0_0_a2_0_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[5]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[5]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[4]_net_1 ), .S(\TM_Packet_Counter_s[5] )
        , .Y(), .FCO(\TM_Packet_Counter_cry[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[14]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[14]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[13]_net_1 ), .S(
        \TM_Packet_Counter_s[14] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[14]_net_1 ));
    SLE \Addr[3]  (.D(\Addr_s[3] ), .CLK(P_CLK), .EN(N_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_USER_RA_TRP1_3));
    CFG4 #( .INIT(16'h0010) )  un1_Flag_B_Tx_Finish17_0_0_o2_RNI47871 
        (.A(Addr), .B(\State[1]_net_1 ), .C(N_1296_i_0), .D(N_1287), 
        .Y(un1_Flag_B_Tx_Finish17_i_0));
    VCC VCC (.Y(VCC_net_1));
    SLE En_ASG (.D(N_29_i_1), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(ENASM));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[16]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[16]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[15]_net_1 ), .S(
        \TM_Packet_Counter_s[16] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[16]_net_1 ));
    SLE \TM_Packet_Counter[20]  (.D(\TM_Packet_Counter_s[20] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[20]));
    SLE \ASM_Count[3]  (.D(N_458_i_0), .CLK(P_CLK), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ASM_Count[3]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \clock_dec_RNI9867[2]  (.A(
        \clock_dec[2]_net_1 ), .B(\clock_dec[1]_net_1 ), .C(
        \clock_dec[0]_net_1 ), .Y(N_1296_i_0));
    CFG4 #( .INIT(16'h777F) )  un1_Flag_B_Tx_Finish17_0_0_o2 (.A(
        pending), .B(En_read_buff), .C(TXD4_net_0), .D(
        Glue_Logic_0_Flag_B_Tx), .Y(N_1287));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[21]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[21]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[20]_net_1 ), .S(
        \TM_Packet_Counter_s[21] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[21]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  USER_REN_TRP1_5_f0_i_0_a2_0 (.A(
        CPU_W_HDL_R_0_USER_RA_TRP1_5), .B(CPU_W_HDL_R_0_USER_RA_TRP1_0)
        , .C(N_1366), .D(N_1346_4), .Y(N_1340));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[6]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[6]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[5]_net_1 ), .S(\TM_Packet_Counter_s[6] )
        , .Y(), .FCO(\TM_Packet_Counter_cry[6]_net_1 ));
    SLE \TM_Packet_Counter[28]  (.D(\TM_Packet_Counter_s[28] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[28]));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_s[31]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[31]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[30]_net_1 ), .S(
        \TM_Packet_Counter_s[31]_net_1 ), .Y(), .FCO());
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[25]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[25]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[24]_net_1 ), .S(
        \TM_Packet_Counter_s[25] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[25]_net_1 ));
    CFG3 #( .INIT(8'h6A) )  \clock_dec_RNO[2]  (.A(
        \clock_dec[2]_net_1 ), .B(\clock_dec[1]_net_1 ), .C(
        \clock_dec[0]_net_1 ), .Y(N_103_i_i_0));
    CFG2 #( .INIT(4'h7) )  \ASM_Count_4_i_0_o3[1]  (.A(
        \ASM_Count[2]_net_1 ), .B(\ASM_Count[3]_net_1 ), .Y(N_1288));
    SLE \Addr[9]  (.D(N_31_i_0), .CLK(P_CLK), .EN(N_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_USER_RA_TRP1_9));
    CFG2 #( .INIT(4'h1) )  \Addr_RNO[9]  (.A(Flag_Type11), .B(
        \State[1]_net_1 ), .Y(N_31_i_0));
    SLE \TM_Packet_Counter[27]  (.D(\TM_Packet_Counter_s[27] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[27]));
    ARI1 #( .INIT(20'h48800) )  \Addr_cry[5]  (.A(VCC_net_1), .B(Addr), 
        .C(CPU_W_HDL_R_0_USER_RA_TRP1_5), .D(GND_net_1), .FCI(
        \Addr_cry[4]_net_1 ), .S(\Addr_s[5] ), .Y(), .FCO(
        \Addr_cry[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[20]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[20]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[19]_net_1 ), .S(
        \TM_Packet_Counter_s[20] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[20]_net_1 ));
    SLE \Addr[0]  (.D(\Addr_s[0] ), .CLK(P_CLK), .EN(N_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_USER_RA_TRP1_0));
    SLE Flag_B_Tx_Finish (.D(Flag_B_Tx_Finish_3), .CLK(P_CLK), .EN(
        N_1296_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CPU_W_HDL_R_0_Flag_B_Tx_Finish));
    CFG2 #( .INIT(4'hE) )  USER_REN_TRP1_5_f0_i_0_o3 (.A(N_1287), .B(
        Addr), .Y(N_1310));
    SLE \TM_Packet_Counter[24]  (.D(\TM_Packet_Counter_s[24] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[24]));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[22]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[22]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[21]_net_1 ), .S(
        \TM_Packet_Counter_s[22] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[22]_net_1 ));
    SLE \TM_Packet_Counter[19]  (.D(\TM_Packet_Counter_s[19] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[19]));
    SLE \TM_Packet_Counter[26]  (.D(\TM_Packet_Counter_s[26] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[26]));
    SLE \TM_Packet_Counter[21]  (.D(\TM_Packet_Counter_s[21] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[21]));
    GND GND (.Y(GND_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[11]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[11]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[10]_net_1 ), .S(
        \TM_Packet_Counter_s[11] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[11]_net_1 ));
    SLE \Addr[4]  (.D(\Addr_s[4] ), .CLK(P_CLK), .EN(N_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_USER_RA_TRP1_4));
    CFG2 #( .INIT(4'h6) )  \clock_dec_RNO[1]  (.A(\clock_dec[0]_net_1 )
        , .B(\clock_dec[1]_net_1 ), .Y(\clock_dec_RNO[1]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \ASM_Count_4_i_0_o3[2]  (.A(
        \ASM_Count[0]_net_1 ), .B(\ASM_Count[1]_net_1 ), .Y(N_85));
    SLE \State[0]  (.D(N_136_i_0), .CLK(P_CLK), .EN(N_1296_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(Addr));
    CFG4 #( .INIT(16'h0045) )  USER_REN_TRP1_RNO (.A(\State[1]_net_1 ), 
        .B(CPU_W_HDL_R_0_USER_REN_TRP1), .C(N_1310), .D(N_1340), .Y(
        N_456_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[15]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[15]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[14]_net_1 ), .S(
        \TM_Packet_Counter_s[15] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[15]_net_1 ));
    SLE \Addr[5]  (.D(\Addr_s[5] ), .CLK(P_CLK), .EN(N_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_USER_RA_TRP1_5));
    SLE \clock_dec[0]  (.D(\clock_dec_i_0[0] ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\clock_dec[0]_net_1 ));
    CFG4 #( .INIT(16'h070F) )  USER_REN_TRP1_5_f0_i_0_a2_0_4_RNIH8LG3 
        (.A(N_1366), .B(CPU_W_HDL_R_0_USER_RA_TRP1_0), .C(
        un1_Flag_B_Tx_Finish17_2_i_i_0_1), .D(N_1346_4), .Y(N_5_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[23]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[23]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[22]_net_1 ), .S(
        \TM_Packet_Counter_s[23] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[23]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[1]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[1]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[0]_net_1 ), .S(\TM_Packet_Counter_s[1] )
        , .Y(), .FCO(\TM_Packet_Counter_cry[1]_net_1 ));
    SLE \TM_Packet_Counter[6]  (.D(\TM_Packet_Counter_s[6] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[6]));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[10]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[10]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[9]_net_1 ), .S(
        \TM_Packet_Counter_s[10] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[10]_net_1 ));
    SLE \TM_Packet_Counter[4]  (.D(\TM_Packet_Counter_s[4] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[4]));
    SLE \TM_Packet_Counter[23]  (.D(\TM_Packet_Counter_s[23] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[23]));
    SLE \TM_Packet_Counter[30]  (.D(\TM_Packet_Counter_s[30] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[30]));
    CFG2 #( .INIT(4'hD) )  Flag_A_Tx_Finish_3_f0_0_0_0_o2 (.A(
        \Flag_Type[0]_net_1 ), .B(\Flag_Type[1]_net_1 ), .Y(N_1292));
    CFG3 #( .INIT(8'h32) )  En_CRC32_RNO (.A(ENCRC), .B(
        \State[1]_net_1 ), .C(Addr), .Y(N_457_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[3]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[3]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[2]_net_1 ), .S(\TM_Packet_Counter_s[3] )
        , .Y(), .FCO(\TM_Packet_Counter_cry[3]_net_1 ));
    SLE \TM_Packet_Counter[10]  (.D(\TM_Packet_Counter_s[10] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[10]));
    SLE \TM_Packet_Counter[3]  (.D(\TM_Packet_Counter_s[3] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[3]));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[0]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[0]), .C(
        GND_net_1), .D(GND_net_1), .FCI(TM_Packet_Counter_cry_cy), .S(
        \TM_Packet_Counter_s[0] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[0]_net_1 ));
    SLE \TM_Packet_Counter[25]  (.D(\TM_Packet_Counter_s[25] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[25]));
    SLE \TM_Packet_Counter[18]  (.D(\TM_Packet_Counter_s[18] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[18]));
    CFG1 #( .INIT(2'h1) )  \clock_dec_RNO[0]  (.A(\clock_dec[0]_net_1 )
        , .Y(\clock_dec_i_0[0] ));
    CFG4 #( .INIT(16'h6E00) )  \ASM_Count_RNO[1]  (.A(
        \ASM_Count[0]_net_1 ), .B(\ASM_Count[1]_net_1 ), .C(N_1288), 
        .D(ENCRC), .Y(N_460_i_0));
    ARI1 #( .INIT(20'h45500) )  \TM_Packet_Counter_cry_cy[0]  (.A(
        VCC_net_1), .B(pos1_En_ASG_net_1), .C(GND_net_1), .D(GND_net_1)
        , .FCI(VCC_net_1), .S(), .Y(), .FCO(TM_Packet_Counter_cry_cy));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[27]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[27]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[26]_net_1 ), .S(
        \TM_Packet_Counter_s[27] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[27]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[12]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[12]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[11]_net_1 ), .S(
        \TM_Packet_Counter_s[12] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[12]_net_1 ));
    SLE \TM_Packet_Counter[17]  (.D(\TM_Packet_Counter_s[17] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[17]));
    SLE \Addr[2]  (.D(\Addr_s[2] ), .CLK(P_CLK), .EN(N_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_USER_RA_TRP1_2));
    SLE \TM_Packet_Counter[8]  (.D(\TM_Packet_Counter_s[8] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[8]));
    SLE \TM_Packet_Counter[22]  (.D(\TM_Packet_Counter_s[22] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[22]));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[7]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[7]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[6]_net_1 ), .S(\TM_Packet_Counter_s[7] )
        , .Y(), .FCO(\TM_Packet_Counter_cry[7]_net_1 ));
    CFG1 #( .INIT(2'h1) )  En_ASG_RNIGT37 (.A(ENASM), .Y(ENASM_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[13]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[13]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[12]_net_1 ), .S(
        \TM_Packet_Counter_s[13] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[13]_net_1 ));
    SLE \State[1]  (.D(\State_ns[1] ), .CLK(P_CLK), .EN(N_1296_i_0), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \State[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  Addr_s_366 (.A(VCC_net_1), .B(Addr), 
        .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), .S(), .Y(), 
        .FCO(Addr_s_366_FCO));
    ARI1 #( .INIT(20'h48800) )  \Addr_cry[4]  (.A(VCC_net_1), .B(Addr), 
        .C(CPU_W_HDL_R_0_USER_RA_TRP1_4), .D(GND_net_1), .FCI(
        \Addr_cry[3]_net_1 ), .S(\Addr_s[4] ), .Y(), .FCO(
        \Addr_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[30]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[30]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[29]_net_1 ), .S(
        \TM_Packet_Counter_s[30] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[30]_net_1 ));
    SLE \TM_Packet_Counter[14]  (.D(\TM_Packet_Counter_s[14] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[14]));
    SLE USER_REN_TRP1 (.D(N_456_i_0), .CLK(P_CLK), .EN(N_1296_i_0), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_USER_REN_TRP1));
    SLE \ASM_Count[2]  (.D(N_459_i_0), .CLK(P_CLK), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ASM_Count[2]_net_1 ));
    CFG4 #( .INIT(16'hFDF5) )  USER_REN_TRP1_5_f0_i_0_a2_1_RNITO242 (
        .A(N_1296_i_0), .B(CPU_W_HDL_R_0_USER_RA_TRP1_5), .C(N_1343), 
        .D(N_1366), .Y(un1_Flag_B_Tx_Finish17_2_i_i_0_1));
    CFG3 #( .INIT(8'h48) )  \ASM_Count_RNO[0]  (.A(
        \ASM_Count[0]_net_1 ), .B(ENCRC), .C(N_1300), .Y(N_461_i_0));
    SLE \TM_Packet_Counter[31]  (.D(\TM_Packet_Counter_s[31]_net_1 ), 
        .CLK(P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[31]));
    SLE \TM_Packet_Counter[16]  (.D(\TM_Packet_Counter_s[16] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[16]));
    ARI1 #( .INIT(20'h48800) )  \Addr_s[7]  (.A(VCC_net_1), .B(Addr), 
        .C(CPU_W_HDL_R_0_USER_RA_TRP1_7), .D(GND_net_1), .FCI(
        \Addr_cry[6]_net_1 ), .S(\Addr_s[7]_net_1 ), .Y(), .FCO());
    CFG3 #( .INIT(8'h04) )  \Addr_RNO_0[9]  (.A(Addr), .B(N_1296_i_0), 
        .C(N_1343), .Y(N_3_i_0));
    SLE \TM_Packet_Counter[11]  (.D(\TM_Packet_Counter_s[11] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[11]));
    SLE \Flag_Type[0]  (.D(Flag_Type11), .CLK(P_CLK), .EN(
        un1_Flag_B_Tx_Finish17_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Flag_Type[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  USER_REN_TRP1_5_f0_i_0_a2_0_4 (.A(
        CPU_W_HDL_R_0_USER_RA_TRP1_4), .B(CPU_W_HDL_R_0_USER_RA_TRP1_3)
        , .C(CPU_W_HDL_R_0_USER_RA_TRP1_2), .D(
        CPU_W_HDL_R_0_USER_RA_TRP1_1), .Y(N_1346_4));
    SLE \TM_Packet_Counter[9]  (.D(\TM_Packet_Counter_s[9] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[9]));
    CFG4 #( .INIT(16'hECA8) )  Flag_B_Tx_Finish_3_f0_0_0_0 (.A(
        \State[1]_net_1 ), .B(CPU_W_HDL_R_0_Flag_B_Tx_Finish), .C(
        Flag_B_Tx_Finish_3_f0_0_0_a2_0_0_net_1), .D(Addr), .Y(
        Flag_B_Tx_Finish_3));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[28]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[28]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[27]_net_1 ), .S(
        \TM_Packet_Counter_s[28] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[28]_net_1 ));
    SLE \ASM_Count[0]  (.D(N_461_i_0), .CLK(P_CLK), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ASM_Count[0]_net_1 ));
    SLE \Addr[7]  (.D(\Addr_s[7]_net_1 ), .CLK(P_CLK), .EN(N_5_i_0), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_USER_RA_TRP1_7));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[17]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[17]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[16]_net_1 ), .S(
        \TM_Packet_Counter_s[17] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[17]_net_1 ));
    CFG4 #( .INIT(16'hAD00) )  \ASM_Count_RNO[2]  (.A(
        \ASM_Count[2]_net_1 ), .B(\ASM_Count[3]_net_1 ), .C(N_85), .D(
        ENCRC), .Y(N_459_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[2]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[2]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[1]_net_1 ), .S(\TM_Packet_Counter_s[2] )
        , .Y(), .FCO(\TM_Packet_Counter_cry[2]_net_1 ));
    SLE En_CRC32 (.D(N_457_i_0), .CLK(P_CLK), .EN(N_1296_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(ENCRC));
    SLE \Flag_Type[1]  (.D(Flag_Type11_i_0), .CLK(P_CLK), .EN(
        un1_Flag_B_Tx_Finish17_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Flag_Type[1]_net_1 ));
    CFG3 #( .INIT(8'h04) )  un1_Flag_B_Tx_Finish17_0_0_o2_RNIRU101 (.A(
        Addr), .B(N_1287), .C(\State[1]_net_1 ), .Y(N_1343));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[29]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[29]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[28]_net_1 ), .S(
        \TM_Packet_Counter_s[29] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[29]_net_1 ));
    SLE \TM_Packet_Counter[7]  (.D(\TM_Packet_Counter_s[7] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[7]));
    SLE \TM_Packet_Counter[13]  (.D(\TM_Packet_Counter_s[13] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[13]));
    ARI1 #( .INIT(20'h48800) )  \Addr_cry[2]  (.A(VCC_net_1), .B(Addr), 
        .C(CPU_W_HDL_R_0_USER_RA_TRP1_2), .D(GND_net_1), .FCI(
        \Addr_cry[1]_net_1 ), .S(\Addr_s[2] ), .Y(), .FCO(
        \Addr_cry[2]_net_1 ));
    CFG4 #( .INIT(16'h0203) )  \State_RNO[0]  (.A(Addr), .B(
        \State[1]_net_1 ), .C(N_1340), .D(N_1287), .Y(N_136_i_0));
    SLE \clock_dec[2]  (.D(N_103_i_i_0), .CLK(P_CLK), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \clock_dec[2]_net_1 ));
    SLE \ASM_Count[1]  (.D(N_460_i_0), .CLK(P_CLK), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \ASM_Count[1]_net_1 ));
    SLE \Addr[1]  (.D(\Addr_s[1] ), .CLK(P_CLK), .EN(N_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_USER_RA_TRP1_1));
    CFG4 #( .INIT(16'hF3A0) )  Flag_A_Tx_Finish_3_f0_0_0_0 (.A(Addr), 
        .B(N_1292), .C(CPU_W_HDL_R_0_Flag_A_Tx_Finish), .D(
        \State[1]_net_1 ), .Y(Flag_A_Tx_Finish_3));
    SLE \TM_Packet_Counter[15]  (.D(\TM_Packet_Counter_s[15] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[15]));
    SLE \TM_Packet_Counter[5]  (.D(\TM_Packet_Counter_s[5] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[5]));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[4]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[4]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[3]_net_1 ), .S(\TM_Packet_Counter_s[4] )
        , .Y(), .FCO(\TM_Packet_Counter_cry[4]_net_1 ));
    SLE \clock_dec[1]  (.D(\clock_dec_RNO[1]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\clock_dec[1]_net_1 ));
    CFG3 #( .INIT(8'h80) )  USER_REN_TRP1_5_f0_i_0_a2_1 (.A(
        CPU_W_HDL_R_0_USER_RA_TRP1_6), .B(Addr), .C(
        CPU_W_HDL_R_0_USER_RA_TRP1_7), .Y(N_1366));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[18]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[18]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[17]_net_1 ), .S(
        \TM_Packet_Counter_s[18] ), .Y(), .FCO(
        \TM_Packet_Counter_cry[18]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  En_ASG_5_i_0_o2 (.A(\ASM_Count[3]_net_1 ), 
        .B(\ASM_Count[1]_net_1 ), .C(\ASM_Count[2]_net_1 ), .Y(N_1300));
    ARI1 #( .INIT(20'h4AA00) )  \TM_Packet_Counter_cry[9]  (.A(
        VCC_net_1), .B(CPU_W_HDL_R_0_TM_Packet_Counter[9]), .C(
        GND_net_1), .D(GND_net_1), .FCI(
        \TM_Packet_Counter_cry[8]_net_1 ), .S(\TM_Packet_Counter_s[9] )
        , .Y(), .FCO(\TM_Packet_Counter_cry[9]_net_1 ));
    SLE \TM_Packet_Counter[12]  (.D(\TM_Packet_Counter_s[12] ), .CLK(
        P_CLK), .EN(ENASM), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CPU_W_HDL_R_0_TM_Packet_Counter[12]));
    
endmodule


module Randomizer(
       pn_reg_0,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       P_CLK,
       S_OUT_0
    );
output pn_reg_0;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  P_CLK;
input  S_OUT_0;

    wire GND_net_1, \pn_reg_3[0]_net_1 , VCC_net_1, \pn_reg[1]_net_1 , 
        \pn_reg_3[1]_net_1 , \pn_reg[2]_net_1 , \pn_reg_3[2]_net_1 , 
        \pn_reg[3]_net_1 , \pn_reg_3[3]_net_1 , \pn_reg[4]_net_1 , 
        \pn_reg_3[4]_net_1 , \pn_reg[5]_net_1 , \pn_reg_3[5]_net_1 , 
        \pn_reg[6]_net_1 , \pn_reg_3[6]_net_1 , \pn_reg[7]_net_1 , 
        \pn_reg_3[7]_net_1 , pn_xorout_0_net_1;
    
    CFG2 #( .INIT(4'hD) )  \pn_reg_3[4]  (.A(S_OUT_0), .B(
        \pn_reg[5]_net_1 ), .Y(\pn_reg_3[4]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \pn_reg_3[1]  (.A(S_OUT_0), .B(
        \pn_reg[2]_net_1 ), .Y(\pn_reg_3[1]_net_1 ));
    SLE \pn_reg[3]  (.D(\pn_reg_3[3]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\pn_reg[3]_net_1 ));
    SLE \pn_reg[0]  (.D(\pn_reg_3[0]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(pn_reg_0));
    SLE \pn_reg[7]  (.D(\pn_reg_3[7]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\pn_reg[7]_net_1 ));
    CFG2 #( .INIT(4'h6) )  pn_xorout_0 (.A(\pn_reg[5]_net_1 ), .B(
        \pn_reg[7]_net_1 ), .Y(pn_xorout_0_net_1));
    SLE \pn_reg[2]  (.D(\pn_reg_3[2]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\pn_reg[2]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'hD) )  \pn_reg_3[5]  (.A(S_OUT_0), .B(
        \pn_reg[6]_net_1 ), .Y(\pn_reg_3[5]_net_1 ));
    SLE \pn_reg[6]  (.D(\pn_reg_3[6]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\pn_reg[6]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \pn_reg_3[3]  (.A(S_OUT_0), .B(
        \pn_reg[4]_net_1 ), .Y(\pn_reg_3[3]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \pn_reg_3[0]  (.A(S_OUT_0), .B(
        \pn_reg[1]_net_1 ), .Y(\pn_reg_3[0]_net_1 ));
    CFG4 #( .INIT(16'h9F6F) )  \pn_reg_3[7]  (.A(\pn_reg[3]_net_1 ), 
        .B(pn_reg_0), .C(S_OUT_0), .D(pn_xorout_0_net_1), .Y(
        \pn_reg_3[7]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \pn_reg_3[6]  (.A(S_OUT_0), .B(
        \pn_reg[7]_net_1 ), .Y(\pn_reg_3[6]_net_1 ));
    SLE \pn_reg[1]  (.D(\pn_reg_3[1]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\pn_reg[1]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \pn_reg_3[2]  (.A(S_OUT_0), .B(
        \pn_reg[3]_net_1 ), .Y(\pn_reg_3[2]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE \pn_reg[4]  (.D(\pn_reg_3[4]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\pn_reg[4]_net_1 ));
    SLE \pn_reg[5]  (.D(\pn_reg_3[5]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\pn_reg[5]_net_1 ));
    
endmodule


module HDL_W_CPU_R_BUFF(
       HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       RX_GPIO1_c,
       EnIP,
       HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish,
       HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish,
       HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1,
       Glue_Logic_0_Flag_B_Rx,
       Flag_RX,
       C_1,
       TC_Decode_0_IP_END_O,
       FALG_FINISH_A_0
    );
output [3:0] HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1;
output [31:0] HDL_W_CPU_R_BUFF_0_MSG_TRP1;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  RX_GPIO1_c;
input  EnIP;
output HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish;
output HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish;
output HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1;
input  Glue_Logic_0_Flag_B_Rx;
input  Flag_RX;
input  C_1;
input  TC_Decode_0_IP_END_O;
input  FALG_FINISH_A_0;

    wire \clk_count[2]_net_1 , VCC_net_1, N_668_i_0, GND_net_1, 
        \clk_count[3]_net_1 , N_667_i_0, \MSG_WA_TRP1_12[0]_net_1 , 
        N_666_i_0, N_665_i_0, \MSG_WA_TRP1_12[3]_net_1 , 
        \Data_A[19]_net_1 , \Data_A_16[19] , 
        Data_A_2_sqmuxa_i_0_0_net_1, \Data_A[20]_net_1 , 
        \Data_A_16[20] , \Data_A[21]_net_1 , \Data_A_16[21] , 
        \Data_A[22]_net_1 , \Data_A_16[22] , \Data_A[23]_net_1 , 
        \Data_A_16[23] , \Data_A[24]_net_1 , \Data_A_16[24] , 
        \Data_A[25]_net_1 , \Data_A_16[25] , \Data_A[26]_net_1 , 
        \Data_A_16[26] , \Data_A[27]_net_1 , \Data_A_16[27] , 
        \Data_A[28]_net_1 , \Data_A_16[28] , \Data_A[29]_net_1 , 
        \Data_A_16[29] , \Data_A[30]_net_1 , \Data_A_16[30] , 
        \Data_A[31]_net_1 , \Data_A_16[31] , \clk_count[0]_net_1 , 
        N_670_i_0, \clk_count[1]_net_1 , N_669_i_0, \Data_A[4]_net_1 , 
        \Data_A_16[4] , \Data_A[5]_net_1 , \Data_A_16[5] , 
        \Data_A[6]_net_1 , \Data_A_16[6] , \Data_A[7]_net_1 , 
        \Data_A_16[7] , \Data_A[8]_net_1 , \Data_A_16[8] , 
        \Data_A[9]_net_1 , \Data_A_16[9] , \Data_A[10]_net_1 , 
        \Data_A_16[10] , \Data_A[11]_net_1 , \Data_A_16[11] , 
        \Data_A[12]_net_1 , \Data_A_16[12] , \Data_A[13]_net_1 , 
        \Data_A_16[13] , \Data_A[14]_net_1 , \Data_A_16[14] , 
        \Data_A[15]_net_1 , \Data_A_16[15] , \Data_A[16]_net_1 , 
        \Data_A_16[16] , \Data_A[17]_net_1 , \Data_A_16[17] , 
        \Data_A[18]_net_1 , \Data_A_16[18] , \Data_B[21]_net_1 , 
        N_1866_i_0, Data_B_0_sqmuxa_i_0_0_net_1, \Data_B[22]_net_1 , 
        N_1849_i_0, \Data_B[23]_net_1 , N_1832_i_0, \Data_B[24]_net_1 , 
        N_1815_i_0, \Data_B[25]_net_1 , N_1798_i_0, \Data_B[26]_net_1 , 
        N_1781_i_0, \Data_B[27]_net_1 , N_1764_i_0, \Data_B[28]_net_1 , 
        N_1747_i_0, \Data_B[29]_net_1 , N_1730_i_0, \Data_B[30]_net_1 , 
        N_1713_i_0, \Data_B[31]_net_1 , N_1696_i_0, \Data_A[0]_net_1 , 
        \Data_A_16[0] , \Data_A[1]_net_1 , \Data_A_16[1] , 
        \Data_A[2]_net_1 , \Data_A_16[2] , \Data_A[3]_net_1 , 
        \Data_A_16[3] , \Data_B[6]_net_1 , N_1679_i_0, 
        \Data_B[7]_net_1 , N_1662_i_0, \Data_B[8]_net_1 , N_1645_i_0, 
        \Data_B[9]_net_1 , N_1628_i_0, \Data_B[10]_net_1 , N_1611_i_0, 
        \Data_B[11]_net_1 , N_1594_i_0, \Data_B[12]_net_1 , N_1577_i_0, 
        \Data_B[13]_net_1 , N_1560_i_0, \Data_B[14]_net_1 , N_1543_i_0, 
        \Data_B[15]_net_1 , N_1526_i_0, \Data_B[16]_net_1 , N_1509_i_0, 
        \Data_B[17]_net_1 , N_1492_i_0, \Data_B[18]_net_1 , N_1475_i_0, 
        \Data_B[19]_net_1 , N_1458_i_0, \Data_B[20]_net_1 , N_1441_i_0, 
        N_1423_i_0, State_Abuff_0_sqmuxa_1_i_o3_0_net_1, N_1403_i_0, 
        N_1383_i_0, N_1363_i_0, N_1343_i_0, N_1323_i_0, N_1303_i_0, 
        N_1283_i_0, N_1263_i_0, \Data_B[0]_net_1 , N_1243_i_0, 
        \Data_B[1]_net_1 , N_1226_i_0, \Data_B[2]_net_1 , N_1209_i_0, 
        \Data_B[3]_net_1 , N_1192_i_0, \Data_B[4]_net_1 , N_1175_i_0, 
        \Data_B[5]_net_1 , N_1158_i_0, N_1140_i_0, N_1120_i_0, 
        N_1100_i_0, N_1080_i_0, N_1060_i_0, N_1040_i_0, N_1020_i_0, 
        N_1000_i_0, N_980_i_0, N_960_i_0, N_940_i_0, N_920_i_0, 
        N_900_i_0, N_880_i_0, N_860_i_0, N_840_i_0, N_820_i_0, 
        N_800_i_0, N_780_i_0, N_760_i_0, N_740_i_0, N_720_i_0, 
        N_700_i_0, Flag_Once_net_1, N_1253, 
        Flag_Once_0_sqmuxa_i_0_0_net_1, Flag_OF_net_1, N_1092_i_0, 
        \State_Abuff[0]_net_1 , State_Abuff_1_sqmuxa, 
        State_Abuff_1_sqmuxa_1_i_0_0_net_1, 
        Flag_A_HDL_Rec_Finish_2_sqmuxa_0_231_a2_0_a2_0_a2_net_1, 
        Flag_A_HDL_Rec_Finish_1_sqmuxa_1_i_0_0_net_1, 
        Flag_B_HDL_Rec_Finish_1_sqmuxa_i_0_0_net_1, N_652_i_0, 
        USER_WEN_TRP1_2_sqmuxa_i_0_0_net_1, \State[0]_net_1 , 
        \State_ns[0] , \State[1]_net_1 , \State_ns[1] , 
        \Bit_Count[0]_net_1 , \Bit_Count_lm[0] , Bit_Counte, 
        \Bit_Count[1]_net_1 , \Bit_Count_lm[1] , \Bit_Count[2]_net_1 , 
        \Bit_Count_lm[2] , \Bit_Count[3]_net_1 , \Bit_Count_lm[3] , 
        \Bit_Count[4]_net_1 , \Bit_Count_lm[4] , \Bit_Count[5]_net_1 , 
        \Bit_Count_lm[5] , \Block_Count[0]_net_1 , \Block_Count_s[0] , 
        Block_Counte, \Block_Count[1]_net_1 , \Block_Count_s[1] , 
        un8lto2, \Block_Count_s[2] , \Block_Count[3]_net_1 , 
        \Block_Count_s[3] , \Block_Count[4]_net_1 , \Block_Count_s[4] , 
        \Block_Count[5]_net_1 , \Block_Count_s[5] , Block_Count_cry_cy, 
        Flag_Once_RNIP8A21_Y, N_159, \Block_Count_cry[0] , 
        \Block_Count_cry[1] , \Block_Count_cry[2] , 
        \Block_Count_cry[3] , \Block_Count_cry[4] , 
        Bit_Count_s_368_FCO, \Bit_Count_cry[1]_net_1 , 
        \Bit_Count_s[1] , \Bit_Count_cry[2]_net_1 , \Bit_Count_s[2] , 
        \Bit_Count_cry[3]_net_1 , \Bit_Count_s[3] , 
        \Bit_Count_s[5]_net_1 , \Bit_Count_cry[4]_net_1 , 
        \Bit_Count_s[4] , N_1097, N_164, N_202_i, N_1108, N_1268, 
        N_1182, \Bit_Count_lm_0_1_0[0]_net_1 , N_500, N_1103, 
        un1_Block_Err_5_0_i_0_net_1, N_1111, N_262_i_0, 
        Data_A_2_sqmuxa_i_0_0_1_net_1, \State_RNIMA5N[0]_net_1 , N_158, 
        \Data_A_16_ns_1[31]_net_1 , Data_A_16_sm0, 
        \Data_A_16_ns_1[30]_net_1 , \Data_A_16_ns_1[29]_net_1 , 
        \Data_A_16_ns_1[28]_net_1 , \Data_A_16_ns_1[27]_net_1 , 
        \Data_A_16_ns_1[26]_net_1 , \Data_A_16_ns_1[25]_net_1 , 
        \Data_A_16_ns_1[24]_net_1 , \Data_A_16_ns_1[23]_net_1 , 
        \Data_A_16_ns_1[22]_net_1 , \Data_A_16_ns_1[21]_net_1 , 
        \Data_A_16_ns_1[20]_net_1 , \Data_A_16_ns_1[19]_net_1 , 
        \Data_A_16_ns_1[18]_net_1 , \Data_A_16_ns_1[17]_net_1 , 
        \Data_A_16_ns_1[16]_net_1 , \Data_A_16_ns_1[15]_net_1 , 
        \Data_A_16_ns_1[14]_net_1 , \Data_A_16_ns_1[13]_net_1 , 
        \Data_A_16_ns_1[12]_net_1 , \Data_A_16_ns_1[11]_net_1 , 
        \Data_A_16_ns_1[10]_net_1 , \Data_A_16_ns_1[9]_net_1 , 
        \Data_A_16_ns_1[8]_net_1 , \Data_A_16_ns_1[7]_net_1 , 
        \Data_A_16_ns_1[6]_net_1 , \Data_A_16_ns_1[5]_net_1 , 
        \Data_A_16_ns_1[4]_net_1 , \Data_A_16_ns_1[3]_net_1 , 
        \Data_A_16_ns_1[2]_net_1 , \Data_A_16_ns_1[1]_net_1 , 
        \Data_A_16_bm[0]_net_1 , \Data_A_16_am[0]_net_1 , N_1275, 
        N_1112, N_1408, N_1124, N_1104, Data_A_1_sqmuxa_sn, 
        Data_B_0_sqmuxa_i_0_0_a2_0_net_1, N_1415, N_290, N_1098, 
        m19_0_0_a2_0, N_1215, N_1257, N_200, \SUM_0[3] , 
        Block_Countlde_0_0_0, un1_Block_Err_3_i_i_o3_0_o2_0, N_1109, 
        \clk_count_6_i_0_1[0]_net_1 , m19_0_0_0, 
        \clk_count_6_i_0_1[2]_net_1 , N_686, 
        MSG_WA_TRP1_0_sqmuxa_1_net_1, N_1255, N_1254, N_1252, N_1114;
    
    SLE \Data_B[8]  (.D(N_1645_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[8]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[22]  (.A(
        \Data_B[22]_net_1 ), .B(\Data_A[22]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_860_i_0));
    SLE \State[0]  (.D(\State_ns[0] ), .CLK(RX_GPIO1_c), .EN(VCC_net_1)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\State[0]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  State_Abuff_1_sqmuxa_1_i_0_0 (.A(N_1112), 
        .B(\State[0]_net_1 ), .C(N_1182), .Y(
        State_Abuff_1_sqmuxa_1_i_0_0_net_1));
    CFG4 #( .INIT(16'h2000) )  MSG_WA_TRP1_0_sqmuxa_1 (.A(EnIP), .B(
        N_1111), .C(\State[0]_net_1 ), .D(
        HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1), .Y(
        MSG_WA_TRP1_0_sqmuxa_1_net_1));
    SLE \MSG_TRP1[21]  (.D(N_880_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[21]));
    SLE \Data_B[2]  (.D(N_1209_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[2]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[8]  (.A(\Data_B[8]_net_1 )
        , .B(\Data_A[8]_net_1 ), .C(N_159), .D(N_158), .Y(N_1140_i_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[16]  (.A(\Data_B[15]_net_1 )
        , .B(\Data_B[16]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1509_i_0));
    CFG4 #( .INIT(16'hECCC) )  \clk_count_6_i_0_a2_RNI274K2[0]  (.A(
        N_1268), .B(un1_Block_Err_3_i_i_o3_0_o2_0), .C(
        TC_Decode_0_IP_END_O), .D(\State[1]_net_1 ), .Y(N_686));
    CFG4 #( .INIT(16'hFFF8) )  \State_RNIAJI01[0]  (.A(
        \State[0]_net_1 ), .B(\State[1]_net_1 ), .C(C_1), .D(
        TC_Decode_0_IP_END_O), .Y(N_1182));
    CFG3 #( .INIT(8'h41) )  \MSG_WA_TRP1_RNO[2]  (.A(N_686), .B(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[2]), .C(N_1114), .Y(N_665_i_0)
        );
    CFG4 #( .INIT(16'h5559) )  \clk_count_6_i_0_x2[3]  (.A(
        \clk_count[3]_net_1 ), .B(\clk_count[0]_net_1 ), .C(N_1097), 
        .D(N_164), .Y(N_202_i));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[10]  (.A(
        \Data_A[9]_net_1 ), .B(\Data_A[10]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[10]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[3]  (.A(
        \Data_A_16_ns_1[3]_net_1 ), .B(\Data_A[3]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[3] ));
    CFG3 #( .INIT(8'h20) )  State_Abuff_1_sqmuxa_0_a3_0_a2 (.A(
        \Bit_Count[5]_net_1 ), .B(\State_Abuff[0]_net_1 ), .C(N_500), 
        .Y(State_Abuff_1_sqmuxa));
    ARI1 #( .INIT(20'h40020) )  Flag_Once_RNIP8A21 (.A(N_159), .B(EnIP)
        , .C(Flag_Once_net_1), .D(\State[0]_net_1 ), .FCI(VCC_net_1), 
        .S(), .Y(Flag_Once_RNIP8A21_Y), .FCO(Block_Count_cry_cy));
    SLE \Data_B[10]  (.D(N_1611_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[10]_net_1 ));
    SLE \Data_A[1]  (.D(\Data_A_16[1] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[1]_net_1 ));
    SLE \Data_B[0]  (.D(N_1243_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[0]_net_1 ));
    SLE \MSG_TRP1[10]  (.D(N_1100_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[10]));
    SLE \Block_Count[3]  (.D(\Block_Count_s[3] ), .CLK(RX_GPIO1_c), 
        .EN(Block_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Block_Count[3]_net_1 ));
    SLE \MSG_TRP1[4]  (.D(N_760_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[4]));
    CFG3 #( .INIT(8'hF8) )  un8lto5_i_a2_0_a2_i_o2 (.A(un8lto2), .B(
        N_1408), .C(N_1415), .Y(N_1111));
    SLE \Data_A[0]  (.D(\Data_A_16[0] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[0]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  \State_ns_1_0_.m22_0_0_a2  (.A(
        \State[0]_net_1 ), .B(EnIP), .C(N_1103), .D(N_159), .Y(N_1252));
    CFG3 #( .INIT(8'h40) )  \Bit_Count_lm_0[4]  (.A(
        \Bit_Count[5]_net_1 ), .B(\Bit_Count_s[4] ), .C(N_500), .Y(
        \Bit_Count_lm[4] ));
    CFG4 #( .INIT(16'hF2F0) )  \State_ns_1_0_.m19_0_0_0  (.A(N_1268), 
        .B(TC_Decode_0_IP_END_O), .C(N_1215), .D(
        Flag_A_HDL_Rec_Finish_2_sqmuxa_0_231_a2_0_a2_0_a2_net_1), .Y(
        m19_0_0_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[20]  (.A(\Data_B[19]_net_1 )
        , .B(\Data_B[20]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1441_i_0));
    SLE \Data_B[5]  (.D(N_1158_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[5]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[12]  (.A(
        \Data_B[12]_net_1 ), .B(\Data_A[12]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1060_i_0));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[24]  (.A(
        \Data_A[23]_net_1 ), .B(\Data_A[24]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[24]_net_1 ));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[23]  (.A(\Data_B[22]_net_1 )
        , .B(\Data_B[23]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1832_i_0));
    SLE \Data_A[6]  (.D(\Data_A_16[6] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[6]_net_1 ));
    CFG4 #( .INIT(16'hF0F8) )  Data_B_0_sqmuxa_i_0_0 (.A(
        Data_B_0_sqmuxa_i_0_0_a2_0_net_1), .B(EnIP), .C(
        \State_RNIMA5N[0]_net_1 ), .D(N_1111), .Y(
        Data_B_0_sqmuxa_i_0_0_net_1));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[31]  (.A(
        \Data_A_16_ns_1[31]_net_1 ), .B(\Data_A[31]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[31] ));
    SLE \MSG_TRP1[20]  (.D(N_900_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[20]));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[4]  (.A(
        \Data_A_16_ns_1[4]_net_1 ), .B(\Data_A[4]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[4] ));
    ARI1 #( .INIT(20'h48800) )  \Block_Count_RNIIM7F2[0]  (.A(
        VCC_net_1), .B(\Block_Count[0]_net_1 ), .C(
        Flag_Once_RNIP8A21_Y), .D(GND_net_1), .FCI(Block_Count_cry_cy), 
        .S(\Block_Count_s[0] ), .Y(), .FCO(\Block_Count_cry[0] ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[22]  (.A(
        \Data_A[21]_net_1 ), .B(\Data_A[22]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[22]_net_1 ));
    SLE \Block_Count[2]  (.D(\Block_Count_s[2] ), .CLK(RX_GPIO1_c), 
        .EN(Block_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(un8lto2));
    SLE \Data_B[14]  (.D(N_1543_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[14]_net_1 ));
    SLE \Data_B[19]  (.D(N_1458_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[19]_net_1 ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[30]  (.A(
        \Data_A[29]_net_1 ), .B(\Data_A[30]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[30]_net_1 ));
    CFG4 #( .INIT(16'hF0F2) )  Flag_OF_RNII5VU1 (.A(N_262_i_0), .B(
        Flag_RX), .C(\State_RNIMA5N[0]_net_1 ), .D(N_1104), .Y(
        un1_Block_Err_3_i_i_o3_0_o2_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_A_16_bm[0]  (.A(\Data_A[0]_net_1 )
        , .B(FALG_FINISH_A_0), .C(\State_RNIMA5N[0]_net_1 ), .D(N_1108)
        , .Y(\Data_A_16_bm[0]_net_1 ));
    SLE \MSG_TRP1[14]  (.D(N_1020_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[14]));
    ARI1 #( .INIT(20'h48800) )  \Block_Count_RNI360M6[3]  (.A(
        VCC_net_1), .B(\Block_Count[3]_net_1 ), .C(
        Flag_Once_RNIP8A21_Y), .D(GND_net_1), .FCI(
        \Block_Count_cry[2] ), .S(\Block_Count_s[3] ), .Y(), .FCO(
        \Block_Count_cry[3] ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[11]  (.A(
        \Data_A_16_ns_1[11]_net_1 ), .B(\Data_A[11]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[11] ));
    CFG4 #( .INIT(16'h020E) )  USER_WEN_TRP1_2_sqmuxa_i_0_0_a2 (.A(
        EnIP), .B(un8lto2), .C(N_1415), .D(N_1408), .Y(N_1275));
    SLE Flag_A_HDL_Rec_Finish (.D(
        Flag_A_HDL_Rec_Finish_2_sqmuxa_0_231_a2_0_a2_0_a2_net_1), .CLK(
        RX_GPIO1_c), .EN(Flag_A_HDL_Rec_Finish_1_sqmuxa_1_i_0_0_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[2]  (.A(\Data_B[1]_net_1 ), 
        .B(\Data_B[2]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 ), 
        .Y(N_1209_i_0));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[22]  (.A(
        \Data_A_16_ns_1[22]_net_1 ), .B(\Data_A[22]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[22] ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[7]  (.A(\Data_B[7]_net_1 )
        , .B(\Data_A[7]_net_1 ), .C(N_159), .D(N_158), .Y(N_700_i_0));
    SLE \MSG_TRP1[16]  (.D(N_980_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[16]));
    SLE \MSG_WA_TRP1[0]  (.D(\MSG_WA_TRP1_12[0]_net_1 ), .CLK(
        RX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0]));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[24]  (.A(
        \Data_B[24]_net_1 ), .B(\Data_A[24]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1403_i_0));
    SLE \MSG_TRP1[12]  (.D(N_1060_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[12]));
    CFG2 #( .INIT(4'h4) )  Flag_Once_RNO (.A(N_159), .B(EnIP), .Y(
        N_1253));
    ARI1 #( .INIT(20'h4AA00) )  \Bit_Count_cry[3]  (.A(VCC_net_1), .B(
        \Bit_Count[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \Bit_Count_cry[2]_net_1 ), .S(\Bit_Count_s[3] ), .Y(), .FCO(
        \Bit_Count_cry[3]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[2]  (.A(
        \Data_A_16_ns_1[2]_net_1 ), .B(\Data_A[2]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[2] ));
    SLE \MSG_TRP1[2]  (.D(N_800_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[2]));
    GND GND (.Y(GND_net_1));
    SLE \Data_B[18]  (.D(N_1475_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[18]_net_1 ));
    CFG4 #( .INIT(16'h3100) )  USER_WEN_TRP1_RNO (.A(EnIP), .B(N_159), 
        .C(\Bit_Count[5]_net_1 ), .D(\State[0]_net_1 ), .Y(N_652_i_0));
    SLE \Bit_Count[5]  (.D(\Bit_Count_lm[5] ), .CLK(RX_GPIO1_c), .EN(
        Bit_Counte), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[5]_net_1 ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[17]  (.A(
        \Data_A[16]_net_1 ), .B(\Data_A[17]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[17]_net_1 ));
    SLE \MSG_TRP1[15]  (.D(N_1000_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[15]));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[25]  (.A(
        \Data_A[24]_net_1 ), .B(\Data_A[25]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[25]_net_1 ));
    CFG4 #( .INIT(16'hAA6A) )  \un1_MSG_WA_TRP1_1.SUM_0[3]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[3]), .B(Flag_RX), .C(N_290), 
        .D(N_1104), .Y(\SUM_0[3] ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[28]  (.A(
        \Data_B[28]_net_1 ), .B(\Data_A[28]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1323_i_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[31]  (.A(\Data_B[30]_net_1 )
        , .B(\Data_B[31]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1696_i_0));
    SLE \Bit_Count[1]  (.D(\Bit_Count_lm[1] ), .CLK(RX_GPIO1_c), .EN(
        Bit_Counte), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[1]_net_1 ));
    SLE \MSG_TRP1[24]  (.D(N_1403_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[24]));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[6]  (.A(
        \Data_A_16_ns_1[6]_net_1 ), .B(\Data_A[6]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[6] ));
    SLE \MSG_WA_TRP1[3]  (.D(\MSG_WA_TRP1_12[3]_net_1 ), .CLK(
        RX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[3]));
    SLE \MSG_TRP1[26]  (.D(N_1363_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[26]));
    SLE \MSG_TRP1[22]  (.D(N_860_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[22]));
    CFG2 #( .INIT(4'h1) )  \State_RNIT3QJ[0]  (.A(\State[1]_net_1 ), 
        .B(\State[0]_net_1 ), .Y(N_262_i_0));
    CFG4 #( .INIT(16'hFDEE) )  \clk_count_6_i_0_1[0]  (.A(
        \clk_count[0]_net_1 ), .B(C_1), .C(TC_Decode_0_IP_END_O), .D(
        N_164), .Y(\clk_count_6_i_0_1[0]_net_1 ));
    CFG4 #( .INIT(16'hDFCC) )  Flag_Once_0_sqmuxa_i_0_0 (.A(EnIP), .B(
        \State_RNIMA5N[0]_net_1 ), .C(Flag_Once_net_1), .D(
        \State[0]_net_1 ), .Y(Flag_Once_0_sqmuxa_i_0_0_net_1));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[7]  (.A(
        \Data_A[6]_net_1 ), .B(\Data_A[7]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[7]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[9]  (.A(
        \Data_A_16_ns_1[9]_net_1 ), .B(\Data_A[9]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[9] ));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[6]  (.A(\Data_B[5]_net_1 ), 
        .B(\Data_B[6]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 ), 
        .Y(N_1679_i_0));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[28]  (.A(
        \Data_A[27]_net_1 ), .B(\Data_A[28]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[28]_net_1 ));
    SLE \Data_A[9]  (.D(\Data_A_16[9] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[9]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[29]  (.A(
        \Data_B[29]_net_1 ), .B(\Data_A[29]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1303_i_0));
    SLE \MSG_TRP1[25]  (.D(N_1383_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[25]));
    CFG2 #( .INIT(4'hE) )  Data_B_12_iv_25_875_i_0_0_o2 (.A(
        \State_Abuff[0]_net_1 ), .B(\Bit_Count[5]_net_1 ), .Y(N_1124));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[11]  (.A(
        \Data_A[10]_net_1 ), .B(\Data_A[11]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[11]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[2]  (.A(\Data_B[2]_net_1 )
        , .B(\Data_A[2]_net_1 ), .C(N_159), .D(N_158), .Y(N_800_i_0));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[14]  (.A(
        \Data_B[14]_net_1 ), .B(\Data_A[14]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1020_i_0));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[20]  (.A(
        \Data_A_16_ns_1[20]_net_1 ), .B(\Data_A[20]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[20] ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[21]  (.A(
        \Data_B[21]_net_1 ), .B(\Data_A[21]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_880_i_0));
    SLE Flag_Once (.D(N_1253), .CLK(RX_GPIO1_c), .EN(
        Flag_Once_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Flag_Once_net_1));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[1]  (.A(\Data_B[0]_net_1 ), 
        .B(\Data_B[1]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 ), 
        .Y(N_1226_i_0));
    SLE \Data_B[15]  (.D(N_1526_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[15]_net_1 ));
    SLE \Data_A[4]  (.D(\Data_A_16[4] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[4]_net_1 ));
    CFG4 #( .INIT(16'h1230) )  \MSG_WA_TRP1_RNO[1]  (.A(
        MSG_WA_TRP1_0_sqmuxa_1_net_1), .B(N_686), .C(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[1]), .D(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0]), .Y(N_666_i_0));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[23]  (.A(
        \Data_A_16_ns_1[23]_net_1 ), .B(\Data_A[23]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[23] ));
    CFG4 #( .INIT(16'hFFDC) )  Data_A_2_sqmuxa_i_0_0 (.A(N_1111), .B(
        N_262_i_0), .C(Data_A_2_sqmuxa_i_0_0_1_net_1), .D(
        \State_RNIMA5N[0]_net_1 ), .Y(Data_A_2_sqmuxa_i_0_0_net_1));
    SLE \MSG_TRP1[31]  (.D(N_1263_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[31]));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[6]  (.A(
        \Data_A[5]_net_1 ), .B(\Data_A[6]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[6]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[30]  (.A(
        \Data_B[30]_net_1 ), .B(\Data_A[30]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1283_i_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[18]  (.A(\Data_B[17]_net_1 )
        , .B(\Data_B[18]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1475_i_0));
    SLE \Block_Count[5]  (.D(\Block_Count_s[5] ), .CLK(RX_GPIO1_c), 
        .EN(Block_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Block_Count[5]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[18]  (.A(
        \Data_B[18]_net_1 ), .B(\Data_A[18]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_940_i_0));
    SLE \Data_B[11]  (.D(N_1594_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[11]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[25]  (.A(
        \Data_A_16_ns_1[25]_net_1 ), .B(\Data_A[25]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[25] ));
    SLE \Block_Count[0]  (.D(\Block_Count_s[0] ), .CLK(RX_GPIO1_c), 
        .EN(Block_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Block_Count[0]_net_1 ));
    CFG4 #( .INIT(16'hF8FF) )  un1_State_4_i_o2 (.A(
        Glue_Logic_0_Flag_B_Rx), .B(Flag_RX), .C(Flag_OF_net_1), .D(
        EnIP), .Y(N_1108));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[3]  (.A(\Data_B[3]_net_1 )
        , .B(\Data_A[3]_net_1 ), .C(N_159), .D(N_158), .Y(N_780_i_0));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[24]  (.A(
        \Data_A_16_ns_1[24]_net_1 ), .B(\Data_A[24]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[24] ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[25]  (.A(
        \Data_B[25]_net_1 ), .B(\Data_A[25]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1383_i_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[26]  (.A(\Data_B[25]_net_1 )
        , .B(\Data_B[26]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1781_i_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[17]  (.A(\Data_B[16]_net_1 )
        , .B(\Data_B[17]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1492_i_0));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[28]  (.A(
        \Data_A_16_ns_1[28]_net_1 ), .B(\Data_A[28]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[28] ));
    SLE \MSG_TRP1[8]  (.D(N_1140_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[8]));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[16]  (.A(
        \Data_A[15]_net_1 ), .B(\Data_A[16]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[16]_net_1 ));
    SLE \Data_B[12]  (.D(N_1577_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[12]_net_1 ));
    SLE \Data_B[17]  (.D(N_1492_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[17]_net_1 ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[9]  (.A(
        \Data_A[8]_net_1 ), .B(\Data_A[9]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[9]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  \un1_MSG_WA_TRP1_1.ANC1_0_o2_i_o2  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[1]), .B(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0]), .C(
        MSG_WA_TRP1_0_sqmuxa_1_net_1), .Y(N_1114));
    ARI1 #( .INIT(20'h48800) )  \Block_Count_RNI0OT28[4]  (.A(
        VCC_net_1), .B(\Block_Count[4]_net_1 ), .C(
        Flag_Once_RNIP8A21_Y), .D(GND_net_1), .FCI(
        \Block_Count_cry[3] ), .S(\Block_Count_s[4] ), .Y(), .FCO(
        \Block_Count_cry[4] ));
    SLE \Block_Count[4]  (.D(\Block_Count_s[4] ), .CLK(RX_GPIO1_c), 
        .EN(Block_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Block_Count[4]_net_1 ));
    SLE \MSG_TRP1[18]  (.D(N_940_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[18]));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[19]  (.A(
        \Data_B[19]_net_1 ), .B(\Data_A[19]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_920_i_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[11]  (.A(\Data_B[10]_net_1 )
        , .B(\Data_B[11]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1594_i_0));
    CFG4 #( .INIT(16'h0103) )  \clk_count_RNO[3]  (.A(N_164), .B(
        N_202_i), .C(C_1), .D(TC_Decode_0_IP_END_O), .Y(N_667_i_0));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[9]  (.A(\Data_B[9]_net_1 )
        , .B(\Data_A[9]_net_1 ), .C(N_159), .D(N_158), .Y(N_1120_i_0));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[31]  (.A(
        \Data_A[30]_net_1 ), .B(\Data_A[31]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[31]_net_1 ));
    CFG3 #( .INIT(8'h40) )  \Bit_Count_lm_0[1]  (.A(
        \Bit_Count[5]_net_1 ), .B(\Bit_Count_s[1] ), .C(N_500), .Y(
        \Bit_Count_lm[1] ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[2]  (.A(
        \Data_A[1]_net_1 ), .B(\Data_A[2]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[2]_net_1 ));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[14]  (.A(\Data_B[13]_net_1 )
        , .B(\Data_B[14]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1543_i_0));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[11]  (.A(
        \Data_B[11]_net_1 ), .B(\Data_A[11]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1080_i_0));
    CFG3 #( .INIT(8'hFB) )  USER_WEN_TRP1_2_sqmuxa_i_0_0 (.A(N_159), 
        .B(\State[0]_net_1 ), .C(N_1275), .Y(
        USER_WEN_TRP1_2_sqmuxa_i_0_0_net_1));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[19]  (.A(
        \Data_A_16_ns_1[19]_net_1 ), .B(\Data_A[19]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[19] ));
    SLE \Data_A[8]  (.D(\Data_A_16[8] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[8]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[17]  (.A(
        \Data_A_16_ns_1[17]_net_1 ), .B(\Data_A[17]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[17] ));
    SLE \MSG_WA_TRP1[1]  (.D(N_666_i_0), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[1]));
    SLE \MSG_TRP1[30]  (.D(N_1283_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[30]));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[29]  (.A(
        \Data_A[28]_net_1 ), .B(\Data_A[29]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[29]_net_1 ));
    SLE \MSG_TRP1[28]  (.D(N_1323_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[28]));
    CFG4 #( .INIT(16'h0302) )  \clk_count_RNO[2]  (.A(N_1097), .B(C_1), 
        .C(\clk_count_6_i_0_1[2]_net_1 ), .D(N_1098), .Y(N_668_i_0));
    SLE \clk_count[0]  (.D(N_670_i_0), .CLK(RX_GPIO1_c), .EN(VCC_net_1)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\clk_count[0]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[15]  (.A(
        \Data_B[15]_net_1 ), .B(\Data_A[15]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1000_i_0));
    CFG3 #( .INIT(8'hBA) )  \State_ns_1_0_.m22_0_0  (.A(N_1252), .B(
        TC_Decode_0_IP_END_O), .C(
        Flag_A_HDL_Rec_Finish_2_sqmuxa_0_231_a2_0_a2_0_a2_net_1), .Y(
        \State_ns[1] ));
    CFG2 #( .INIT(4'h1) )  \Data_A_16_am_RNO[0]  (.A(
        \State_Abuff[0]_net_1 ), .B(\State[1]_net_1 ), .Y(
        Data_A_1_sqmuxa_sn));
    SLE \MSG_TRP1[7]  (.D(N_700_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[7]));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[8]  (.A(\Data_B[7]_net_1 ), 
        .B(\Data_B[8]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 ), 
        .Y(N_1645_i_0));
    SLE \Data_B[16]  (.D(N_1509_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[16]_net_1 ));
    CFG4 #( .INIT(16'hBB0F) )  \Bit_Count_lm_0[0]  (.A(
        \Bit_Count[5]_net_1 ), .B(\Bit_Count[0]_net_1 ), .C(
        \Bit_Count_lm_0_1_0[0]_net_1 ), .D(N_500), .Y(
        \Bit_Count_lm[0] ));
    SLE \Data_B[1]  (.D(N_1226_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \Bit_Count_cry[4]  (.A(VCC_net_1), .B(
        \Bit_Count[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \Bit_Count_cry[3]_net_1 ), .S(\Bit_Count_s[4] ), .Y(), .FCO(
        \Bit_Count_cry[4]_net_1 ));
    CFG3 #( .INIT(8'h01) )  un1_Block_Err_5_0_i_a2_0 (.A(N_159), .B(
        \State[0]_net_1 ), .C(N_1108), .Y(N_1215));
    SLE \Data_A[10]  (.D(\Data_A_16[10] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[10]_net_1 ));
    SLE \Data_A[5]  (.D(\Data_A_16[5] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[5]_net_1 ));
    SLE \MSG_TRP1[5]  (.D(N_740_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[5]));
    SLE \Data_A[20]  (.D(\Data_A_16[20] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[20]_net_1 ));
    SLE \Data_B[13]  (.D(N_1560_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[13]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[16]  (.A(
        \Data_A_16_ns_1[16]_net_1 ), .B(\Data_A[16]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[16] ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[14]  (.A(
        \Data_A[13]_net_1 ), .B(\Data_A[14]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[14]_net_1 ));
    SLE \Bit_Count[4]  (.D(\Bit_Count_lm[4] ), .CLK(RX_GPIO1_c), .EN(
        Bit_Counte), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[4]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \clk_count_6_i_0_o2_0[2]  (.A(
        \clk_count[1]_net_1 ), .B(\clk_count[2]_net_1 ), .Y(N_1097));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[5]  (.A(
        \Data_A_16_ns_1[5]_net_1 ), .B(\Data_A[5]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[5] ));
    ARI1 #( .INIT(20'h4AA00) )  \Bit_Count_cry[1]  (.A(VCC_net_1), .B(
        \Bit_Count[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        Bit_Count_s_368_FCO), .S(\Bit_Count_s[1] ), .Y(), .FCO(
        \Bit_Count_cry[1]_net_1 ));
    SLE \MSG_TRP1[17]  (.D(N_960_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[17]));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[19]  (.A(\Data_B[18]_net_1 )
        , .B(\Data_B[19]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1458_i_0));
    CFG3 #( .INIT(8'h12) )  \MSG_WA_TRP1_12[0]  (.A(
        MSG_WA_TRP1_0_sqmuxa_1_net_1), .B(N_686), .C(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0]), .Y(
        \MSG_WA_TRP1_12[0]_net_1 ));
    CFG4 #( .INIT(16'h3B00) )  Data_A_2_sqmuxa_i_0_0_1 (.A(EnIP), .B(
        N_158), .C(\Bit_Count[5]_net_1 ), .D(\State[0]_net_1 ), .Y(
        Data_A_2_sqmuxa_i_0_0_1_net_1));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[5]  (.A(\Data_B[5]_net_1 )
        , .B(\Data_A[5]_net_1 ), .C(N_159), .D(N_158), .Y(N_740_i_0));
    CFG2 #( .INIT(4'hD) )  Flag_OF_RNI5IHI (.A(EnIP), .B(Flag_OF_net_1)
        , .Y(N_1104));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[12]  (.A(
        \Data_A[11]_net_1 ), .B(\Data_A[12]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[12]_net_1 ));
    SLE \Data_B[9]  (.D(N_1628_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[9]_net_1 ));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[15]  (.A(\Data_B[14]_net_1 )
        , .B(\Data_B[15]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1526_i_0));
    SLE \Data_B[20]  (.D(N_1441_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[20]_net_1 ));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[5]  (.A(\Data_B[4]_net_1 ), 
        .B(\Data_B[5]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 ), 
        .Y(N_1158_i_0));
    SLE \Data_A[2]  (.D(\Data_A_16[2] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[2]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[8]  (.A(
        \Data_A_16_ns_1[8]_net_1 ), .B(\Data_A[8]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[8] ));
    CFG2 #( .INIT(4'h1) )  
        Flag_A_HDL_Rec_Finish_2_sqmuxa_0_231_a2_0_a2_0_a2 (.A(N_164), 
        .B(C_1), .Y(
        Flag_A_HDL_Rec_Finish_2_sqmuxa_0_231_a2_0_a2_0_a2_net_1));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[4]  (.A(
        \Data_A[3]_net_1 ), .B(\Data_A[4]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[4]_net_1 ));
    SLE \Data_A[14]  (.D(\Data_A_16[14] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[14]_net_1 ));
    SLE \clk_count[2]  (.D(N_668_i_0), .CLK(RX_GPIO1_c), .EN(VCC_net_1)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\clk_count[2]_net_1 ));
    SLE \Data_A[7]  (.D(\Data_A_16[7] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[7]_net_1 ));
    SLE \Data_A[19]  (.D(\Data_A_16[19] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[19]_net_1 ));
    SLE \Data_A[24]  (.D(\Data_A_16[24] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[24]_net_1 ));
    CFG4 #( .INIT(16'hCD01) )  \clk_count_6_i_0_o2[1]  (.A(N_1097), .B(
        N_164), .C(\clk_count[3]_net_1 ), .D(TC_Decode_0_IP_END_O), .Y(
        N_1109));
    SLE \MSG_TRP1[27]  (.D(N_1343_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[27]));
    SLE \Data_A[29]  (.D(\Data_A_16[29] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[29]_net_1 ));
    SLE \Data_B[3]  (.D(N_1192_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[3]_net_1 ));
    CFG4 #( .INIT(16'hFFF4) )  Flag_A_HDL_Rec_Finish_1_sqmuxa_1_i_0_0 
        (.A(Flag_RX), .B(N_262_i_0), .C(\State_RNIMA5N[0]_net_1 ), .D(
        N_1254), .Y(Flag_A_HDL_Rec_Finish_1_sqmuxa_1_i_0_0_net_1));
    CFG3 #( .INIT(8'h10) )  \State_ns_1_0_.m19_0_0_a2_0_0  (.A(N_159), 
        .B(TC_Decode_0_IP_END_O), .C(\State[0]_net_1 ), .Y(
        m19_0_0_a2_0));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[23]  (.A(
        \Data_A[22]_net_1 ), .B(\Data_A[23]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[23]_net_1 ));
    SLE \MSG_TRP1[9]  (.D(N_1120_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[9]));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[15]  (.A(
        \Data_A[14]_net_1 ), .B(\Data_A[15]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[15]_net_1 ));
    SLE \Data_A[30]  (.D(\Data_A_16[30] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[30]_net_1 ));
    SLE \Data_A[18]  (.D(\Data_A_16[18] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[18]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[4]  (.A(\Data_B[4]_net_1 )
        , .B(\Data_A[4]_net_1 ), .C(N_159), .D(N_158), .Y(N_760_i_0));
    SLE Flag_B_HDL_Rec_Finish (.D(
        Flag_A_HDL_Rec_Finish_2_sqmuxa_0_231_a2_0_a2_0_a2_net_1), .CLK(
        RX_GPIO1_c), .EN(Flag_B_HDL_Rec_Finish_1_sqmuxa_i_0_0_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish));
    SLE \Data_B[4]  (.D(N_1175_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[4]_net_1 ));
    CFG4 #( .INIT(16'hF3F1) )  \clk_count_6_i_0_1[2]  (.A(
        \clk_count[1]_net_1 ), .B(\clk_count[2]_net_1 ), .C(N_1109), 
        .D(N_1098), .Y(\clk_count_6_i_0_1[2]_net_1 ));
    CFG4 #( .INIT(16'h00FB) )  \Bit_Count_lm_0_1_0[0]  (.A(
        TC_Decode_0_IP_END_O), .B(N_1103), .C(N_159), .D(
        un1_Block_Err_5_0_i_0_net_1), .Y(\Bit_Count_lm_0_1_0[0]_net_1 )
        );
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[21]  (.A(
        \Data_A_16_ns_1[21]_net_1 ), .B(\Data_A[21]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[21] ));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[30]  (.A(\Data_B[29]_net_1 )
        , .B(\Data_B[30]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1713_i_0));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[23]  (.A(
        \Data_B[23]_net_1 ), .B(\Data_A[23]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1423_i_0));
    CFG3 #( .INIT(8'h4C) )  Data_B_0_sqmuxa_i_0_0_a2_0 (.A(
        \Bit_Count[5]_net_1 ), .B(\State[0]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .Y(Data_B_0_sqmuxa_i_0_0_a2_0_net_1));
    SLE \Data_B[24]  (.D(N_1815_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[24]_net_1 ));
    SLE \Data_A[28]  (.D(\Data_A_16[28] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[28]_net_1 ));
    SLE \Data_B[29]  (.D(N_1730_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[29]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  \Data_A_16_ns[0]  (.A(
        \Data_A_16_bm[0]_net_1 ), .B(Data_A_16_sm0), .C(
        \Data_A_16_am[0]_net_1 ), .Y(\Data_A_16[0] ));
    SLE \Data_B[6]  (.D(N_1679_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[6]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[1]  (.A(\Data_B[1]_net_1 )
        , .B(\Data_A[1]_net_1 ), .C(N_159), .D(N_158), .Y(N_820_i_0));
    SLE \MSG_TRP1[1]  (.D(N_820_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[1]));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[28]  (.A(\Data_B[27]_net_1 )
        , .B(\Data_B[28]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1747_i_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[12]  (.A(\Data_B[11]_net_1 )
        , .B(\Data_B[12]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1577_i_0));
    CFG2 #( .INIT(4'h7) )  Data_A_2_sqmuxa_i_0_0_o2 (.A(EnIP), .B(
        \State_Abuff[0]_net_1 ), .Y(N_158));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[18]  (.A(
        \Data_A[17]_net_1 ), .B(\Data_A[18]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[18]_net_1 ));
    SLE \clk_count[1]  (.D(N_669_i_0), .CLK(RX_GPIO1_c), .EN(VCC_net_1)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\clk_count[1]_net_1 ));
    SLE \Data_B[7]  (.D(N_1662_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[7]_net_1 ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[20]  (.A(
        \Data_A[19]_net_1 ), .B(\Data_A[20]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[20]_net_1 ));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[27]  (.A(\Data_B[26]_net_1 )
        , .B(\Data_B[27]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1764_i_0));
    SLE \Data_B[30]  (.D(N_1713_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[30]_net_1 ));
    SLE \Data_B[28]  (.D(N_1747_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[28]_net_1 ));
    CFG2 #( .INIT(4'hB) )  \clk_count_6_i_0_o2[0]  (.A(N_164), .B(
        \clk_count[0]_net_1 ), .Y(N_1098));
    CFG4 #( .INIT(16'h00C6) )  \MSG_WA_TRP1_12[3]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[2]), .B(\SUM_0[3] ), .C(
        N_1114), .D(N_686), .Y(\MSG_WA_TRP1_12[3]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[1]  (.A(
        \Data_A_16_ns_1[1]_net_1 ), .B(\Data_A[1]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[1] ));
    CFG4 #( .INIT(16'h2000) )  Flag_B_HDL_Rec_Finish_1_sqmuxa_i_0_0_a2 
        (.A(N_1268), .B(N_200), .C(TC_Decode_0_IP_END_O), .D(
        \State[1]_net_1 ), .Y(N_1255));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[21]  (.A(\Data_B[20]_net_1 )
        , .B(\Data_B[21]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1866_i_0));
    ARI1 #( .INIT(20'h4AA00) )  Bit_Count_s_368 (.A(VCC_net_1), .B(
        \Bit_Count[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(Bit_Count_s_368_FCO));
    SLE \Bit_Count[0]  (.D(\Bit_Count_lm[0] ), .CLK(RX_GPIO1_c), .EN(
        Bit_Counte), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[0]_net_1 ));
    SLE \Data_A[15]  (.D(\Data_A_16[15] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[15]_net_1 ));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[24]  (.A(\Data_B[23]_net_1 )
        , .B(\Data_B[24]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1815_i_0));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[13]  (.A(
        \Data_B[13]_net_1 ), .B(\Data_A[13]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1040_i_0));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[12]  (.A(
        \Data_A_16_ns_1[12]_net_1 ), .B(\Data_A[12]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[12] ));
    SLE \Data_A[25]  (.D(\Data_A_16[25] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[25]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[27]  (.A(
        \Data_B[27]_net_1 ), .B(\Data_A[27]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1343_i_0));
    CFG4 #( .INIT(16'hCECC) )  Flag_Once_RNID7HP1 (.A(EnIP), .B(N_1182)
        , .C(Flag_Once_net_1), .D(\State[0]_net_1 ), .Y(
        Block_Countlde_0_0_0));
    SLE \Data_A[11]  (.D(\Data_A_16[11] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[11]_net_1 ));
    CFG3 #( .INIT(8'h40) )  \Bit_Count_lm_0[2]  (.A(
        \Bit_Count[5]_net_1 ), .B(\Bit_Count_s[2] ), .C(N_500), .Y(
        \Bit_Count_lm[2] ));
    CFG2 #( .INIT(4'hE) )  MSG_TRP1_11_iv_28_304_i_0_0_o2 (.A(
        \State[1]_net_1 ), .B(C_1), .Y(N_159));
    SLE \MSG_TRP1[13]  (.D(N_1040_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[13]));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[4]  (.A(\Data_B[3]_net_1 ), 
        .B(\Data_B[4]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 ), 
        .Y(N_1175_i_0));
    SLE \Data_A[21]  (.D(\Data_A_16[21] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[21]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[0]  (.A(\Data_B[0]_net_1 )
        , .B(\Data_A[0]_net_1 ), .C(N_159), .D(N_158), .Y(N_840_i_0));
    SLE \MSG_TRP1[3]  (.D(N_780_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[3]));
    SLE \Data_A[12]  (.D(\Data_A_16[12] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[12]_net_1 ));
    SLE \Data_A[17]  (.D(\Data_A_16[17] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[17]_net_1 ));
    CFG4 #( .INIT(16'hAAAC) )  \Data_A_16_am[0]  (.A(FALG_FINISH_A_0), 
        .B(\Data_A[0]_net_1 ), .C(\Bit_Count[5]_net_1 ), .D(
        Data_A_1_sqmuxa_sn), .Y(\Data_A_16_am[0]_net_1 ));
    CFG2 #( .INIT(4'h2) )  Flag_B_HDL_Rec_Finish_1_sqmuxa_i_0_0_a2_0 (
        .A(N_262_i_0), .B(Glue_Logic_0_Flag_B_Rx), .Y(N_290));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[10]  (.A(\Data_B[9]_net_1 ), 
        .B(\Data_B[10]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 ), 
        .Y(N_1611_i_0));
    CFG4 #( .INIT(16'hFEFA) )  
        USER_WEN_TRP1_2_sqmuxa_i_0_0_a2_RNI38L42 (.A(N_1182), .B(
        \State[0]_net_1 ), .C(N_1257), .D(N_1275), .Y(Bit_Counte));
    CFG2 #( .INIT(4'hE) )  Data_A_16s2 (.A(\State_RNIMA5N[0]_net_1 ), 
        .B(N_262_i_0), .Y(Data_A_16_sm0));
    SLE \State[1]  (.D(\State_ns[1] ), .CLK(RX_GPIO1_c), .EN(VCC_net_1)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\State[1]_net_1 ));
    SLE \Data_B[25]  (.D(N_1798_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[25]_net_1 ));
    CFG4 #( .INIT(16'hCCCD) )  un1_Block_Err_5_0_i_0 (.A(
        \State[0]_net_1 ), .B(N_1215), .C(C_1), .D(
        TC_Decode_0_IP_END_O), .Y(un1_Block_Err_5_0_i_0_net_1));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[20]  (.A(
        \Data_B[20]_net_1 ), .B(\Data_A[20]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_900_i_0));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[26]  (.A(
        \Data_B[26]_net_1 ), .B(\Data_A[26]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1363_i_0));
    SLE \Data_A[22]  (.D(\Data_A_16[22] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[22]_net_1 ));
    SLE \Data_A[27]  (.D(\Data_A_16[27] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[27]_net_1 ));
    SLE \MSG_TRP1[0]  (.D(N_840_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[0]));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[6]  (.A(\Data_B[6]_net_1 )
        , .B(\Data_A[6]_net_1 ), .C(N_159), .D(N_158), .Y(N_720_i_0));
    CFG4 #( .INIT(16'h0401) )  \clk_count_RNO[1]  (.A(C_1), .B(
        \clk_count[1]_net_1 ), .C(N_1109), .D(N_1098), .Y(N_669_i_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[13]  (.A(\Data_B[12]_net_1 )
        , .B(\Data_B[13]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1560_i_0));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[30]  (.A(
        \Data_A_16_ns_1[30]_net_1 ), .B(\Data_A[30]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[30] ));
    SLE \MSG_TRP1[23]  (.D(N_1423_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[23]));
    SLE \Data_B[21]  (.D(N_1866_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[21]_net_1 ));
    CFG3 #( .INIT(8'hC4) )  State_Abuff_0_sqmuxa_1_i_o3_0_o2 (.A(EnIP), 
        .B(N_1275), .C(\Bit_Count[5]_net_1 ), .Y(N_1112));
    CFG3 #( .INIT(8'hFE) )  Flag_B_HDL_Rec_Finish_1_sqmuxa_i_0_0 (.A(
        N_1255), .B(N_290), .C(\State_RNIMA5N[0]_net_1 ), .Y(
        Flag_B_HDL_Rec_Finish_1_sqmuxa_i_0_0_net_1));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[19]  (.A(
        \Data_A[18]_net_1 ), .B(\Data_A[19]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[19]_net_1 ));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[7]  (.A(\Data_B[6]_net_1 ), 
        .B(\Data_B[7]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 ), 
        .Y(N_1662_i_0));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[27]  (.A(
        \Data_A[26]_net_1 ), .B(\Data_A[27]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[27]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \clk_count_6_i_0_o2[3]  (.A(
        \State[1]_net_1 ), .B(\State[0]_net_1 ), .Y(N_164));
    SLE \clk_count[3]  (.D(N_667_i_0), .CLK(RX_GPIO1_c), .EN(VCC_net_1)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\clk_count[3]_net_1 ));
    CFG3 #( .INIT(8'hEC) )  State_Abuff_0_sqmuxa_1_i_o3_0 (.A(
        \State[0]_net_1 ), .B(\State_RNIMA5N[0]_net_1 ), .C(N_1112), 
        .Y(State_Abuff_0_sqmuxa_1_i_o3_0_net_1));
    CFG3 #( .INIT(8'hEA) )  \State_RNIMA5N[0]  (.A(C_1), .B(
        \State[0]_net_1 ), .C(\State[1]_net_1 ), .Y(
        \State_RNIMA5N[0]_net_1 ));
    SLE \Bit_Count[2]  (.D(\Bit_Count_lm[2] ), .CLK(RX_GPIO1_c), .EN(
        Bit_Counte), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[2]_net_1 ));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[3]  (.A(\Data_B[2]_net_1 ), 
        .B(\Data_B[3]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 ), 
        .Y(N_1192_i_0));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[29]  (.A(\Data_B[28]_net_1 )
        , .B(\Data_B[29]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1730_i_0));
    SLE \Data_B[22]  (.D(N_1849_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[22]_net_1 ));
    SLE \Data_B[27]  (.D(N_1764_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[27]_net_1 ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[17]  (.A(
        \Data_B[17]_net_1 ), .B(\Data_A[17]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_960_i_0));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[31]  (.A(
        \Data_B[31]_net_1 ), .B(\Data_A[31]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1263_i_0));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[10]  (.A(
        \Data_A_16_ns_1[10]_net_1 ), .B(\Data_A[10]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[10] ));
    CFG3 #( .INIT(8'hFE) )  un8lto5_i_a2_0_a2_i_o2_0 (.A(
        \Block_Count[5]_net_1 ), .B(\Block_Count[4]_net_1 ), .C(
        \Block_Count[3]_net_1 ), .Y(N_1415));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[5]  (.A(
        \Data_A[4]_net_1 ), .B(\Data_A[5]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[5]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[7]  (.A(
        \Data_A_16_ns_1[7]_net_1 ), .B(\Data_A[7]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[7] ));
    SLE \MSG_TRP1[19]  (.D(N_920_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[19]));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[25]  (.A(\Data_B[24]_net_1 )
        , .B(\Data_B[25]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1798_i_0));
    SLE \Data_A[16]  (.D(\Data_A_16[16] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[16]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[29]  (.A(
        \Data_A_16_ns_1[29]_net_1 ), .B(\Data_A[29]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[29] ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[13]  (.A(
        \Data_A_16_ns_1[13]_net_1 ), .B(\Data_A[13]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[13] ));
    CFG2 #( .INIT(4'h1) )  \clk_count_RNO[0]  (.A(
        \clk_count_6_i_0_1[0]_net_1 ), .B(N_1268), .Y(N_670_i_0));
    SLE \MSG_TRP1[6]  (.D(N_720_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[6]));
    SLE \Data_A[31]  (.D(\Data_A_16[31] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[31]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \Block_Count_RNO[5]  (.A(VCC_net_1), 
        .B(\Block_Count[5]_net_1 ), .C(Flag_Once_RNIP8A21_Y), .D(
        GND_net_1), .FCI(\Block_Count_cry[4] ), .S(\Block_Count_s[5] ), 
        .Y(), .FCO());
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[27]  (.A(
        \Data_A_16_ns_1[27]_net_1 ), .B(\Data_A[27]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[27] ));
    ARI1 #( .INIT(20'h4AA00) )  \Bit_Count_cry[2]  (.A(VCC_net_1), .B(
        \Bit_Count[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \Bit_Count_cry[1]_net_1 ), .S(\Bit_Count_s[2] ), .Y(), .FCO(
        \Bit_Count_cry[2]_net_1 ));
    CFG4 #( .INIT(16'hFF02) )  un1_Block_Err_5_0_i_o2_RNI33K72 (.A(
        \State[0]_net_1 ), .B(EnIP), .C(N_1103), .D(
        Block_Countlde_0_0_0), .Y(Block_Counte));
    SLE \Data_A[26]  (.D(\Data_A_16[26] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[26]_net_1 ));
    SLE \Data_A[3]  (.D(\Data_A_16[3] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[3]_net_1 ));
    SLE \MSG_WA_TRP1[2]  (.D(N_665_i_0), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[2]));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[15]  (.A(
        \Data_A_16_ns_1[15]_net_1 ), .B(\Data_A[15]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[15] ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[10]  (.A(
        \Data_B[10]_net_1 ), .B(\Data_A[10]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_1100_i_0));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[14]  (.A(
        \Data_A_16_ns_1[14]_net_1 ), .B(\Data_A[14]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[14] ));
    CFG4 #( .INIT(16'h0C0A) )  \MSG_TRP1_RNO[16]  (.A(
        \Data_B[16]_net_1 ), .B(\Data_A[16]_net_1 ), .C(N_159), .D(
        N_158), .Y(N_980_i_0));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[21]  (.A(
        \Data_A[20]_net_1 ), .B(\Data_A[21]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[21]_net_1 ));
    SLE \Data_A[13]  (.D(\Data_A_16[13] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[13]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[18]  (.A(
        \Data_A_16_ns_1[18]_net_1 ), .B(\Data_A[18]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[18] ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[1]  (.A(
        \Data_A[0]_net_1 ), .B(\Data_A[1]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[1]_net_1 ));
    CFG3 #( .INIT(8'hFD) )  un1_Block_Err_5_0_i_o2 (.A(un8lto2), .B(
        N_1408), .C(N_1415), .Y(N_1103));
    CFG2 #( .INIT(4'hE) )  \State_ns_1_0_.m19_0_o2_4_i_o2  (.A(
        \Block_Count[0]_net_1 ), .B(\Block_Count[1]_net_1 ), .Y(N_1408)
        );
    ARI1 #( .INIT(20'h48800) )  \Block_Count_RNIC55S3[1]  (.A(
        VCC_net_1), .B(\Block_Count[1]_net_1 ), .C(
        Flag_Once_RNIP8A21_Y), .D(GND_net_1), .FCI(
        \Block_Count_cry[0] ), .S(\Block_Count_s[1] ), .Y(), .FCO(
        \Block_Count_cry[1] ));
    SLE \Block_Count[1]  (.D(\Block_Count_s[1] ), .CLK(RX_GPIO1_c), 
        .EN(Block_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Block_Count[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  un1_State_4_i_o2_RNIHKCO (.A(N_1108), .B(
        N_262_i_0), .Y(N_1257));
    CFG4 #( .INIT(16'hEEEC) )  \State_ns_1_0_.m19_0_0  (.A(
        m19_0_0_a2_0), .B(m19_0_0_0), .C(EnIP), .D(N_1103), .Y(
        \State_ns[0] ));
    SLE \MSG_TRP1[29]  (.D(N_1303_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[29]));
    SLE \Data_A[23]  (.D(\Data_A_16[23] ), .CLK(RX_GPIO1_c), .EN(
        Data_A_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_A[23]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  
        Flag_A_HDL_Rec_Finish_1_sqmuxa_1_i_0_0_a2 (.A(N_1268), .B(
        N_200), .C(TC_Decode_0_IP_END_O), .D(\State[1]_net_1 ), .Y(
        N_1254));
    CFG4 #( .INIT(16'h0020) )  \clk_count_6_i_0_a2[0]  (.A(
        \clk_count[2]_net_1 ), .B(\clk_count[3]_net_1 ), .C(
        \clk_count[1]_net_1 ), .D(\clk_count[0]_net_1 ), .Y(N_1268));
    SLE \Bit_Count[3]  (.D(\Bit_Count_lm[3] ), .CLK(RX_GPIO1_c), .EN(
        Bit_Counte), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[3]_net_1 ));
    SLE USER_WEN_TRP1 (.D(N_652_i_0), .CLK(RX_GPIO1_c), .EN(
        USER_WEN_TRP1_2_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1));
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[9]  (.A(\Data_B[8]_net_1 ), 
        .B(\Data_B[9]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 ), 
        .Y(N_1628_i_0));
    SLE \Data_B[26]  (.D(N_1781_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[26]_net_1 ));
    SLE \Data_B[31]  (.D(N_1696_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[31]_net_1 ));
    CFG3 #( .INIT(8'h40) )  \Bit_Count_lm_0[5]  (.A(
        \Bit_Count[5]_net_1 ), .B(\Bit_Count_s[5]_net_1 ), .C(N_500), 
        .Y(\Bit_Count_lm[5] ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[8]  (.A(
        \Data_A[7]_net_1 ), .B(\Data_A[8]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[8]_net_1 ));
    CFG4 #( .INIT(16'h06C6) )  \Data_A_16_ns[26]  (.A(
        \Data_A_16_ns_1[26]_net_1 ), .B(\Data_A[26]_net_1 ), .C(
        Data_A_16_sm0), .D(\State_RNIMA5N[0]_net_1 ), .Y(
        \Data_A_16[26] ));
    SLE \State_Abuff[0]  (.D(State_Abuff_1_sqmuxa), .CLK(RX_GPIO1_c), 
        .EN(State_Abuff_1_sqmuxa_1_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \State_Abuff[0]_net_1 ));
    CFG4 #( .INIT(16'h00CA) )  \Data_B_RNO[0]  (.A(\Data_B[0]_net_1 ), 
        .B(FALG_FINISH_A_0), .C(N_1124), .D(N_159), .Y(N_1243_i_0));
    SLE Flag_OF (.D(EnIP), .CLK(RX_GPIO1_c), .EN(N_1092_i_0), .ALn(
        VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), 
        .LAT(GND_net_1), .Q(Flag_OF_net_1));
    CFG4 #( .INIT(16'h0020) )  Flag_OF_RNO (.A(N_1108), .B(N_159), .C(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .D(\State[0]_net_1 )
        , .Y(N_1092_i_0));
    SLE \MSG_TRP1[11]  (.D(N_1080_i_0), .CLK(RX_GPIO1_c), .EN(
        State_Abuff_0_sqmuxa_1_i_o3_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[11]));
    CFG4 #( .INIT(16'h5557) )  
        Flag_A_HDL_Rec_Finish_1_sqmuxa_1_i_0_0_o2 (.A(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[3]), .B(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[2]), .C(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[1]), .D(
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0]), .Y(N_200));
    ARI1 #( .INIT(20'h48800) )  \Block_Count_RNI7L295[2]  (.A(
        VCC_net_1), .B(Flag_Once_RNIP8A21_Y), .C(un8lto2), .D(
        GND_net_1), .FCI(\Block_Count_cry[1] ), .S(\Block_Count_s[2] ), 
        .Y(), .FCO(\Block_Count_cry[2] ));
    SLE \Data_B[23]  (.D(N_1832_i_0), .CLK(RX_GPIO1_c), .EN(
        Data_B_0_sqmuxa_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_B[23]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \Bit_Count_s[5]  (.A(VCC_net_1), .B(
        \Bit_Count[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \Bit_Count_cry[4]_net_1 ), .S(\Bit_Count_s[5]_net_1 ), .Y(), 
        .FCO());
    CFG4 #( .INIT(16'h0A0C) )  \Data_B_RNO[22]  (.A(\Data_B[21]_net_1 )
        , .B(\Data_B[22]_net_1 ), .C(N_159), .D(\State_Abuff[0]_net_1 )
        , .Y(N_1849_i_0));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[3]  (.A(
        \Data_A[2]_net_1 ), .B(\Data_A[3]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[3]_net_1 ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[26]  (.A(
        \Data_A[25]_net_1 ), .B(\Data_A[26]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[26]_net_1 ));
    CFG4 #( .INIT(16'h0006) )  \Data_A_16_ns_1[13]  (.A(
        \Data_A[12]_net_1 ), .B(\Data_A[13]_net_1 ), .C(
        \State_Abuff[0]_net_1 ), .D(\State[1]_net_1 ), .Y(
        \Data_A_16_ns_1[13]_net_1 ));
    CFG4 #( .INIT(16'h0008) )  un1_Block_Err_5_0_i_a2_2 (.A(
        \State[0]_net_1 ), .B(EnIP), .C(N_1111), .D(N_159), .Y(N_500));
    CFG3 #( .INIT(8'h40) )  \Bit_Count_lm_0[3]  (.A(
        \Bit_Count[5]_net_1 ), .B(\Bit_Count_s[3] ), .C(N_500), .Y(
        \Bit_Count_lm[3] ));
    
endmodule


module DATA_OUT(
       shift1_reg_4,
       shift1_reg_0,
       TX_GPIO0_c,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       TX_GPIO1_c,
       Convolutional_Encoder_out_1_0,
       P_CLK
    );
input  shift1_reg_4;
input  shift1_reg_0;
output TX_GPIO0_c;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  TX_GPIO1_c;
input  Convolutional_Encoder_out_1_0;
input  P_CLK;

    wire VCC_net_1, DataO_2_net_1, GND_net_1;
    
    CFG4 #( .INIT(16'h65A9) )  DataO_2 (.A(
        Convolutional_Encoder_out_1_0), .B(P_CLK), .C(shift1_reg_4), 
        .D(shift1_reg_0), .Y(DataO_2_net_1));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    SLE DataO (.D(DataO_2_net_1), .CLK(TX_GPIO1_c), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TX_GPIO0_c));
    
endmodule


module COREAPB3_MUXPTOB3(
       CoreAPB3_0_APBmslave3_PRDATA,
       test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA,
       test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx,
       iPSELS_raw23,
       CoreAPB3_0_APBmslave3_PREADY,
       N_623_i_0
    );
input  [31:0] CoreAPB3_0_APBmslave3_PRDATA;
output [31:0] test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA;
input  test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx;
input  iPSELS_raw23;
input  CoreAPB3_0_APBmslave3_PREADY;
output N_623_i_0;

    wire GND_net_1, VCC_net_1;
    
    CFG3 #( .INIT(8'h80) )  \PRDATA[29]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[29]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[29]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[14]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[14]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[14]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[4]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[4]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[4]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[25]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[25]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[25]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[10]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[10]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[10]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[2]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[2]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[2]));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h80) )  \PRDATA[31]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[31]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[31]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[1]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[1]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[1]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[8]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[8]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[8]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[12]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[12]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[12]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[27]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[27]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[27]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[19]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[19]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[19]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[23]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[23]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[23]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[5]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[5]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[5]));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h80) )  \PRDATA[26]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[26]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[26]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[30]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[30]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[30]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[15]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[15]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[15]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[0]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[0]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[0]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[3]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[3]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[3]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[28]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[28]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[28]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[21]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[21]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[21]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[17]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[17]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[17]));
    CFG3 #( .INIT(8'hF7) )  N_623_i (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PREADY), .Y(N_623_i_0));
    CFG3 #( .INIT(8'h80) )  \PRDATA[24]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[24]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[24]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[9]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[9]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[9]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[6]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[6]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[6]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[13]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[13]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[13]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[16]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[16]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[16]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[20]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[20]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[20]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[7]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[7]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[7]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[18]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[18]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[18]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[11]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[11]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[11]));
    CFG3 #( .INIT(8'h80) )  \PRDATA[22]  (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        iPSELS_raw23), .C(CoreAPB3_0_APBmslave3_PRDATA[22]), .Y(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[22]));
    
endmodule


module CoreAPB3_Z1(
       CoreAPB3_0_APBmslave3_PADDR,
       CoreAPB3_0_APBmslave3_PRDATA,
       test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA,
       iPSELS_raw23,
       test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx,
       CoreAPB3_0_APBmslave3_PREADY,
       N_623_i_0
    );
input  [31:28] CoreAPB3_0_APBmslave3_PADDR;
input  [31:0] CoreAPB3_0_APBmslave3_PRDATA;
output [31:0] test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA;
output iPSELS_raw23;
input  test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx;
input  CoreAPB3_0_APBmslave3_PREADY;
output N_623_i_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    COREAPB3_MUXPTOB3 u_mux_p_to_b3 (.CoreAPB3_0_APBmslave3_PRDATA({
        CoreAPB3_0_APBmslave3_PRDATA[31], 
        CoreAPB3_0_APBmslave3_PRDATA[30], 
        CoreAPB3_0_APBmslave3_PRDATA[29], 
        CoreAPB3_0_APBmslave3_PRDATA[28], 
        CoreAPB3_0_APBmslave3_PRDATA[27], 
        CoreAPB3_0_APBmslave3_PRDATA[26], 
        CoreAPB3_0_APBmslave3_PRDATA[25], 
        CoreAPB3_0_APBmslave3_PRDATA[24], 
        CoreAPB3_0_APBmslave3_PRDATA[23], 
        CoreAPB3_0_APBmslave3_PRDATA[22], 
        CoreAPB3_0_APBmslave3_PRDATA[21], 
        CoreAPB3_0_APBmslave3_PRDATA[20], 
        CoreAPB3_0_APBmslave3_PRDATA[19], 
        CoreAPB3_0_APBmslave3_PRDATA[18], 
        CoreAPB3_0_APBmslave3_PRDATA[17], 
        CoreAPB3_0_APBmslave3_PRDATA[16], 
        CoreAPB3_0_APBmslave3_PRDATA[15], 
        CoreAPB3_0_APBmslave3_PRDATA[14], 
        CoreAPB3_0_APBmslave3_PRDATA[13], 
        CoreAPB3_0_APBmslave3_PRDATA[12], 
        CoreAPB3_0_APBmslave3_PRDATA[11], 
        CoreAPB3_0_APBmslave3_PRDATA[10], 
        CoreAPB3_0_APBmslave3_PRDATA[9], 
        CoreAPB3_0_APBmslave3_PRDATA[8], 
        CoreAPB3_0_APBmslave3_PRDATA[7], 
        CoreAPB3_0_APBmslave3_PRDATA[6], 
        CoreAPB3_0_APBmslave3_PRDATA[5], 
        CoreAPB3_0_APBmslave3_PRDATA[4], 
        CoreAPB3_0_APBmslave3_PRDATA[3], 
        CoreAPB3_0_APBmslave3_PRDATA[2], 
        CoreAPB3_0_APBmslave3_PRDATA[1], 
        CoreAPB3_0_APBmslave3_PRDATA[0]}), 
        .test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA({
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[31], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[30], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[29], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[28], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[27], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[26], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[25], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[24], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[23], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[22], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[21], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[20], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[19], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[18], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[17], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[16], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[15], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[14], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[13], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[12], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[11], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[10], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[9], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[8], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[7], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[6], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[5], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[4], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[3], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[2], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[1], 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[0]}), 
        .test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), 
        .iPSELS_raw23(iPSELS_raw23), .CoreAPB3_0_APBmslave3_PREADY(
        CoreAPB3_0_APBmslave3_PREADY), .N_623_i_0(N_623_i_0));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h0400) )  iPSELS_raw23_inst_1 (.A(
        CoreAPB3_0_APBmslave3_PADDR[31]), .B(
        CoreAPB3_0_APBmslave3_PADDR[28]), .C(
        CoreAPB3_0_APBmslave3_PADDR[30]), .D(
        CoreAPB3_0_APBmslave3_PADDR[29]), .Y(iPSELS_raw23));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_18(
       synd_w,
       CODE_FROM_RAM_27,
       CODE_FROM_RAM_24,
       CODE_FROM_RAM_22,
       CODE_FROM_RAM_28,
       CODE_FROM_RAM_35,
       CODE_FROM_RAM_14,
       CODE_FROM_RAM_10,
       CODE_FROM_RAM_8,
       CODE_FROM_RAM_13,
       CODE_FROM_RAM_5,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_17,
       CODE_FROM_RAM_19,
       CODE_FROM_RAM_34,
       CODE_FROM_RAM_31
    );
output [2:2] synd_w;
input  CODE_FROM_RAM_27;
input  CODE_FROM_RAM_24;
input  CODE_FROM_RAM_22;
input  CODE_FROM_RAM_28;
input  CODE_FROM_RAM_35;
input  CODE_FROM_RAM_14;
input  CODE_FROM_RAM_10;
input  CODE_FROM_RAM_8;
input  CODE_FROM_RAM_13;
input  CODE_FROM_RAM_5;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_17;
input  CODE_FROM_RAM_19;
input  CODE_FROM_RAM_34;
input  CODE_FROM_RAM_31;

    wire \outp_9[0]_net_1 , \outp_3[0]_net_1 , \outp_2[0] , 
        \outp_8[0]_net_1 , GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_3[0]  (.A(CODE_FROM_RAM_35), .B(
        CODE_FROM_RAM_14), .C(CODE_FROM_RAM_10), .D(CODE_FROM_RAM_8), 
        .Y(\outp_3[0]_net_1 ));
    CFG3 #( .INIT(8'h96) )  \outp_2_0[0]  (.A(CODE_FROM_RAM_13), .B(
        CODE_FROM_RAM_5), .C(CODE_FROM_RAM_0), .Y(\outp_2[0] ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(CODE_FROM_RAM_34), .B(
        CODE_FROM_RAM_31), .C(\outp_9[0]_net_1 ), .D(\outp_8[0]_net_1 )
        , .Y(synd_w[2]));
    CFG4 #( .INIT(16'h6996) )  \outp_9[0]  (.A(CODE_FROM_RAM_27), .B(
        CODE_FROM_RAM_24), .C(CODE_FROM_RAM_22), .D(CODE_FROM_RAM_28), 
        .Y(\outp_9[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp_8[0]  (.A(\outp_3[0]_net_1 ), .B(
        \outp_2[0] ), .C(CODE_FROM_RAM_17), .D(CODE_FROM_RAM_19), .Y(
        \outp_8[0]_net_1 ));
    
endmodule


module wide_xor_15s_3s_4294967295_4294967295_3s_4_1(
       synd_w,
       CODE_FROM_RAM_27,
       CODE_FROM_RAM_24,
       CODE_FROM_RAM_22,
       CODE_FROM_RAM_28,
       CODE_FROM_RAM_35,
       CODE_FROM_RAM_14,
       CODE_FROM_RAM_10,
       CODE_FROM_RAM_8,
       CODE_FROM_RAM_13,
       CODE_FROM_RAM_5,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_17,
       CODE_FROM_RAM_19,
       CODE_FROM_RAM_34,
       CODE_FROM_RAM_31
    );
output [2:2] synd_w;
input  CODE_FROM_RAM_27;
input  CODE_FROM_RAM_24;
input  CODE_FROM_RAM_22;
input  CODE_FROM_RAM_28;
input  CODE_FROM_RAM_35;
input  CODE_FROM_RAM_14;
input  CODE_FROM_RAM_10;
input  CODE_FROM_RAM_8;
input  CODE_FROM_RAM_13;
input  CODE_FROM_RAM_5;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_17;
input  CODE_FROM_RAM_19;
input  CODE_FROM_RAM_34;
input  CODE_FROM_RAM_31;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_18 \genXOR[2].layer_xor_0  (.synd_w({
        synd_w[2]}), .CODE_FROM_RAM_27(CODE_FROM_RAM_27), 
        .CODE_FROM_RAM_24(CODE_FROM_RAM_24), .CODE_FROM_RAM_22(
        CODE_FROM_RAM_22), .CODE_FROM_RAM_28(CODE_FROM_RAM_28), 
        .CODE_FROM_RAM_35(CODE_FROM_RAM_35), .CODE_FROM_RAM_14(
        CODE_FROM_RAM_14), .CODE_FROM_RAM_10(CODE_FROM_RAM_10), 
        .CODE_FROM_RAM_8(CODE_FROM_RAM_8), .CODE_FROM_RAM_13(
        CODE_FROM_RAM_13), .CODE_FROM_RAM_5(CODE_FROM_RAM_5), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM_0), .CODE_FROM_RAM_17(
        CODE_FROM_RAM_17), .CODE_FROM_RAM_19(CODE_FROM_RAM_19), 
        .CODE_FROM_RAM_34(CODE_FROM_RAM_34), .CODE_FROM_RAM_31(
        CODE_FROM_RAM_31));
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_16(
       synd_w,
       CODE_FROM_RAM_34,
       CODE_FROM_RAM_33,
       CODE_FROM_RAM_30,
       CODE_FROM_RAM_28,
       CODE_FROM_RAM_38,
       CODE_FROM_RAM_16,
       CODE_FROM_RAM_14,
       CODE_FROM_RAM_9,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_7,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_25,
       CODE_FROM_RAM_23,
       CODE_FROM_RAM_19,
       CODE_FROM_RAM_20
    );
output [0:0] synd_w;
input  CODE_FROM_RAM_34;
input  CODE_FROM_RAM_33;
input  CODE_FROM_RAM_30;
input  CODE_FROM_RAM_28;
input  CODE_FROM_RAM_38;
input  CODE_FROM_RAM_16;
input  CODE_FROM_RAM_14;
input  CODE_FROM_RAM_9;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_7;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_25;
input  CODE_FROM_RAM_23;
input  CODE_FROM_RAM_19;
input  CODE_FROM_RAM_20;

    wire \outp_11[0]_net_1 , \outp_4[0]_net_1 , \outp_5[0]_net_1 , 
        \outp_10[0]_net_1 , GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h6996) )  \outp_4[0]  (.A(CODE_FROM_RAM_38), .B(
        CODE_FROM_RAM_16), .C(CODE_FROM_RAM_14), .D(CODE_FROM_RAM_9), 
        .Y(\outp_4[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_5[0]  (.A(\outp_4[0]_net_1 ), .B(
        CODE_FROM_RAM_11), .C(CODE_FROM_RAM_7), .D(CODE_FROM_RAM_0), 
        .Y(\outp_5[0]_net_1 ));
    CFG3 #( .INIT(8'h96) )  \outp_10[0]  (.A(\outp_5[0]_net_1 ), .B(
        CODE_FROM_RAM_25), .C(CODE_FROM_RAM_23), .Y(\outp_10[0]_net_1 )
        );
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(CODE_FROM_RAM_19), .B(
        CODE_FROM_RAM_20), .C(\outp_11[0]_net_1 ), .D(
        \outp_10[0]_net_1 ), .Y(synd_w[0]));
    CFG4 #( .INIT(16'h6996) )  \outp_11[0]  (.A(CODE_FROM_RAM_34), .B(
        CODE_FROM_RAM_33), .C(CODE_FROM_RAM_30), .D(CODE_FROM_RAM_28), 
        .Y(\outp_11[0]_net_1 ));
    
endmodule


module wide_xor_15s_3s_4294967295_4294967295_3s_4(
       synd_w,
       CODE_FROM_RAM_34,
       CODE_FROM_RAM_33,
       CODE_FROM_RAM_30,
       CODE_FROM_RAM_28,
       CODE_FROM_RAM_38,
       CODE_FROM_RAM_16,
       CODE_FROM_RAM_14,
       CODE_FROM_RAM_9,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_7,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_25,
       CODE_FROM_RAM_23,
       CODE_FROM_RAM_19,
       CODE_FROM_RAM_20
    );
output [0:0] synd_w;
input  CODE_FROM_RAM_34;
input  CODE_FROM_RAM_33;
input  CODE_FROM_RAM_30;
input  CODE_FROM_RAM_28;
input  CODE_FROM_RAM_38;
input  CODE_FROM_RAM_16;
input  CODE_FROM_RAM_14;
input  CODE_FROM_RAM_9;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_7;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_25;
input  CODE_FROM_RAM_23;
input  CODE_FROM_RAM_19;
input  CODE_FROM_RAM_20;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_16 \genXOR[2].layer_xor_0  (.synd_w({
        synd_w[0]}), .CODE_FROM_RAM_34(CODE_FROM_RAM_34), 
        .CODE_FROM_RAM_33(CODE_FROM_RAM_33), .CODE_FROM_RAM_30(
        CODE_FROM_RAM_30), .CODE_FROM_RAM_28(CODE_FROM_RAM_28), 
        .CODE_FROM_RAM_38(CODE_FROM_RAM_38), .CODE_FROM_RAM_16(
        CODE_FROM_RAM_16), .CODE_FROM_RAM_14(CODE_FROM_RAM_14), 
        .CODE_FROM_RAM_9(CODE_FROM_RAM_9), .CODE_FROM_RAM_11(
        CODE_FROM_RAM_11), .CODE_FROM_RAM_7(CODE_FROM_RAM_7), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM_0), .CODE_FROM_RAM_25(
        CODE_FROM_RAM_25), .CODE_FROM_RAM_23(CODE_FROM_RAM_23), 
        .CODE_FROM_RAM_19(CODE_FROM_RAM_19), .CODE_FROM_RAM_20(
        CODE_FROM_RAM_20));
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_21(
       synd_w_5,
       synd_w,
       CODE_FROM_RAM_26,
       CODE_FROM_RAM_25,
       CODE_FROM_RAM_18,
       CODE_FROM_RAM_15,
       CODE_FROM_RAM_32,
       CODE_FROM_RAM_10,
       CODE_FROM_RAM_3,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_8,
       CODE_FROM_RAM_6,
       CODE_FROM_RAM_13,
       CODE_FROM_RAM_29
    );
input  [5:5] synd_w_5;
output [5:5] synd_w;
input  CODE_FROM_RAM_26;
input  CODE_FROM_RAM_25;
input  CODE_FROM_RAM_18;
input  CODE_FROM_RAM_15;
input  CODE_FROM_RAM_32;
input  CODE_FROM_RAM_10;
input  CODE_FROM_RAM_3;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_8;
input  CODE_FROM_RAM_6;
input  CODE_FROM_RAM_13;
input  CODE_FROM_RAM_29;

    wire \outp_8[0]_net_1 , \outp_2[0] , \outp_4[0]_net_1 , GND_net_1, 
        VCC_net_1;
    
    CFG4 #( .INIT(16'h6996) )  \outp_4[0]  (.A(CODE_FROM_RAM_8), .B(
        CODE_FROM_RAM_6), .C(\outp_2[0] ), .D(CODE_FROM_RAM_13), .Y(
        \outp_4[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_2_0[0]  (.A(CODE_FROM_RAM_32), .B(
        CODE_FROM_RAM_10), .C(CODE_FROM_RAM_3), .D(CODE_FROM_RAM_0), 
        .Y(\outp_2[0] ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(synd_w_5[5]), .B(
        CODE_FROM_RAM_29), .C(\outp_4[0]_net_1 ), .D(\outp_8[0]_net_1 )
        , .Y(synd_w[5]));
    CFG4 #( .INIT(16'h6996) )  \outp_8[0]  (.A(CODE_FROM_RAM_26), .B(
        CODE_FROM_RAM_25), .C(CODE_FROM_RAM_18), .D(CODE_FROM_RAM_15), 
        .Y(\outp_8[0]_net_1 ));
    
endmodule


module wide_xor_15s_3s_4294967295_4294967295_3s_4_4(
       synd_w_5,
       synd_w,
       CODE_FROM_RAM_26,
       CODE_FROM_RAM_25,
       CODE_FROM_RAM_18,
       CODE_FROM_RAM_15,
       CODE_FROM_RAM_32,
       CODE_FROM_RAM_10,
       CODE_FROM_RAM_3,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_8,
       CODE_FROM_RAM_6,
       CODE_FROM_RAM_13,
       CODE_FROM_RAM_29
    );
input  [5:5] synd_w_5;
output [5:5] synd_w;
input  CODE_FROM_RAM_26;
input  CODE_FROM_RAM_25;
input  CODE_FROM_RAM_18;
input  CODE_FROM_RAM_15;
input  CODE_FROM_RAM_32;
input  CODE_FROM_RAM_10;
input  CODE_FROM_RAM_3;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_8;
input  CODE_FROM_RAM_6;
input  CODE_FROM_RAM_13;
input  CODE_FROM_RAM_29;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_21 \genXOR[2].layer_xor_0  (.synd_w_5({
        synd_w_5[5]}), .synd_w({synd_w[5]}), .CODE_FROM_RAM_26(
        CODE_FROM_RAM_26), .CODE_FROM_RAM_25(CODE_FROM_RAM_25), 
        .CODE_FROM_RAM_18(CODE_FROM_RAM_18), .CODE_FROM_RAM_15(
        CODE_FROM_RAM_15), .CODE_FROM_RAM_32(CODE_FROM_RAM_32), 
        .CODE_FROM_RAM_10(CODE_FROM_RAM_10), .CODE_FROM_RAM_3(
        CODE_FROM_RAM_3), .CODE_FROM_RAM_0(CODE_FROM_RAM_0), 
        .CODE_FROM_RAM_8(CODE_FROM_RAM_8), .CODE_FROM_RAM_6(
        CODE_FROM_RAM_6), .CODE_FROM_RAM_13(CODE_FROM_RAM_13), 
        .CODE_FROM_RAM_29(CODE_FROM_RAM_29));
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_20(
       synd_w,
       CODE_FROM_RAM_28,
       CODE_FROM_RAM_24,
       CODE_FROM_RAM_22,
       CODE_FROM_RAM_21,
       CODE_FROM_RAM_34,
       CODE_FROM_RAM_13,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_9,
       CODE_FROM_RAM_6,
       CODE_FROM_RAM_4,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_16,
       CODE_FROM_RAM_18,
       CODE_FROM_RAM_32,
       CODE_FROM_RAM_29
    );
output [4:4] synd_w;
input  CODE_FROM_RAM_28;
input  CODE_FROM_RAM_24;
input  CODE_FROM_RAM_22;
input  CODE_FROM_RAM_21;
input  CODE_FROM_RAM_34;
input  CODE_FROM_RAM_13;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_9;
input  CODE_FROM_RAM_6;
input  CODE_FROM_RAM_4;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_16;
input  CODE_FROM_RAM_18;
input  CODE_FROM_RAM_32;
input  CODE_FROM_RAM_29;

    wire \outp_10[0]_net_1 , \outp_4[0]_net_1 , \outp_3[0]_net_1 , 
        \outp_9[0]_net_1 , GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h6996) )  \outp_4[0]  (.A(CODE_FROM_RAM_34), .B(
        CODE_FROM_RAM_13), .C(CODE_FROM_RAM_11), .D(CODE_FROM_RAM_9), 
        .Y(\outp_4[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h96) )  \outp_3[0]  (.A(CODE_FROM_RAM_6), .B(
        CODE_FROM_RAM_4), .C(CODE_FROM_RAM_0), .Y(\outp_3[0]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_10[0]  (.A(CODE_FROM_RAM_28), .B(
        CODE_FROM_RAM_24), .C(CODE_FROM_RAM_22), .D(CODE_FROM_RAM_21), 
        .Y(\outp_10[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(CODE_FROM_RAM_32), .B(
        CODE_FROM_RAM_29), .C(\outp_10[0]_net_1 ), .D(
        \outp_9[0]_net_1 ), .Y(synd_w[4]));
    CFG4 #( .INIT(16'h6996) )  \outp_9[0]  (.A(\outp_4[0]_net_1 ), .B(
        \outp_3[0]_net_1 ), .C(CODE_FROM_RAM_16), .D(CODE_FROM_RAM_18), 
        .Y(\outp_9[0]_net_1 ));
    
endmodule


module wide_xor_15s_3s_4294967295_4294967295_3s_4_3(
       synd_w,
       CODE_FROM_RAM_28,
       CODE_FROM_RAM_24,
       CODE_FROM_RAM_22,
       CODE_FROM_RAM_21,
       CODE_FROM_RAM_34,
       CODE_FROM_RAM_13,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_9,
       CODE_FROM_RAM_6,
       CODE_FROM_RAM_4,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_16,
       CODE_FROM_RAM_18,
       CODE_FROM_RAM_32,
       CODE_FROM_RAM_29
    );
output [4:4] synd_w;
input  CODE_FROM_RAM_28;
input  CODE_FROM_RAM_24;
input  CODE_FROM_RAM_22;
input  CODE_FROM_RAM_21;
input  CODE_FROM_RAM_34;
input  CODE_FROM_RAM_13;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_9;
input  CODE_FROM_RAM_6;
input  CODE_FROM_RAM_4;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_16;
input  CODE_FROM_RAM_18;
input  CODE_FROM_RAM_32;
input  CODE_FROM_RAM_29;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_20 \genXOR[2].layer_xor_0  (.synd_w({
        synd_w[4]}), .CODE_FROM_RAM_28(CODE_FROM_RAM_28), 
        .CODE_FROM_RAM_24(CODE_FROM_RAM_24), .CODE_FROM_RAM_22(
        CODE_FROM_RAM_22), .CODE_FROM_RAM_21(CODE_FROM_RAM_21), 
        .CODE_FROM_RAM_34(CODE_FROM_RAM_34), .CODE_FROM_RAM_13(
        CODE_FROM_RAM_13), .CODE_FROM_RAM_11(CODE_FROM_RAM_11), 
        .CODE_FROM_RAM_9(CODE_FROM_RAM_9), .CODE_FROM_RAM_6(
        CODE_FROM_RAM_6), .CODE_FROM_RAM_4(CODE_FROM_RAM_4), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM_0), .CODE_FROM_RAM_16(
        CODE_FROM_RAM_16), .CODE_FROM_RAM_18(CODE_FROM_RAM_18), 
        .CODE_FROM_RAM_32(CODE_FROM_RAM_32), .CODE_FROM_RAM_29(
        CODE_FROM_RAM_29));
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_17(
       synd_w,
       CODE_FROM_RAM_34,
       CODE_FROM_RAM_31,
       CODE_FROM_RAM_30,
       CODE_FROM_RAM_27,
       CODE_FROM_RAM_36,
       CODE_FROM_RAM_16,
       CODE_FROM_RAM_13,
       CODE_FROM_RAM_8,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_6,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_22,
       CODE_FROM_RAM_25,
       CODE_FROM_RAM_20,
       CODE_FROM_RAM_17
    );
output [1:1] synd_w;
input  CODE_FROM_RAM_34;
input  CODE_FROM_RAM_31;
input  CODE_FROM_RAM_30;
input  CODE_FROM_RAM_27;
input  CODE_FROM_RAM_36;
input  CODE_FROM_RAM_16;
input  CODE_FROM_RAM_13;
input  CODE_FROM_RAM_8;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_6;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_22;
input  CODE_FROM_RAM_25;
input  CODE_FROM_RAM_20;
input  CODE_FROM_RAM_17;

    wire \outp_10[0]_net_1 , \outp_3[0] , \outp_2[0]_net_1 , 
        \outp_9[0]_net_1 , GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_3_0[0]  (.A(CODE_FROM_RAM_36), .B(
        CODE_FROM_RAM_16), .C(CODE_FROM_RAM_13), .D(CODE_FROM_RAM_8), 
        .Y(\outp_3[0] ));
    CFG3 #( .INIT(8'h96) )  \outp_2[0]  (.A(CODE_FROM_RAM_11), .B(
        CODE_FROM_RAM_6), .C(CODE_FROM_RAM_0), .Y(\outp_2[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp_10[0]  (.A(CODE_FROM_RAM_34), .B(
        CODE_FROM_RAM_31), .C(CODE_FROM_RAM_30), .D(CODE_FROM_RAM_27), 
        .Y(\outp_10[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(CODE_FROM_RAM_20), .B(
        CODE_FROM_RAM_17), .C(\outp_10[0]_net_1 ), .D(
        \outp_9[0]_net_1 ), .Y(synd_w[1]));
    CFG4 #( .INIT(16'h6996) )  \outp_9[0]  (.A(\outp_3[0] ), .B(
        \outp_2[0]_net_1 ), .C(CODE_FROM_RAM_22), .D(CODE_FROM_RAM_25), 
        .Y(\outp_9[0]_net_1 ));
    
endmodule


module wide_xor_15s_3s_4294967295_4294967295_3s_4_0(
       synd_w,
       CODE_FROM_RAM_34,
       CODE_FROM_RAM_31,
       CODE_FROM_RAM_30,
       CODE_FROM_RAM_27,
       CODE_FROM_RAM_36,
       CODE_FROM_RAM_16,
       CODE_FROM_RAM_13,
       CODE_FROM_RAM_8,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_6,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_22,
       CODE_FROM_RAM_25,
       CODE_FROM_RAM_20,
       CODE_FROM_RAM_17
    );
output [1:1] synd_w;
input  CODE_FROM_RAM_34;
input  CODE_FROM_RAM_31;
input  CODE_FROM_RAM_30;
input  CODE_FROM_RAM_27;
input  CODE_FROM_RAM_36;
input  CODE_FROM_RAM_16;
input  CODE_FROM_RAM_13;
input  CODE_FROM_RAM_8;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_6;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_22;
input  CODE_FROM_RAM_25;
input  CODE_FROM_RAM_20;
input  CODE_FROM_RAM_17;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_17 \genXOR[2].layer_xor_0  (.synd_w({
        synd_w[1]}), .CODE_FROM_RAM_34(CODE_FROM_RAM_34), 
        .CODE_FROM_RAM_31(CODE_FROM_RAM_31), .CODE_FROM_RAM_30(
        CODE_FROM_RAM_30), .CODE_FROM_RAM_27(CODE_FROM_RAM_27), 
        .CODE_FROM_RAM_36(CODE_FROM_RAM_36), .CODE_FROM_RAM_16(
        CODE_FROM_RAM_16), .CODE_FROM_RAM_13(CODE_FROM_RAM_13), 
        .CODE_FROM_RAM_8(CODE_FROM_RAM_8), .CODE_FROM_RAM_11(
        CODE_FROM_RAM_11), .CODE_FROM_RAM_6(CODE_FROM_RAM_6), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM_0), .CODE_FROM_RAM_22(
        CODE_FROM_RAM_22), .CODE_FROM_RAM_25(CODE_FROM_RAM_25), 
        .CODE_FROM_RAM_20(CODE_FROM_RAM_20), .CODE_FROM_RAM_17(
        CODE_FROM_RAM_17));
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_19(
       synd_w_5,
       synd_w,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_5,
       CODE_FROM_RAM_21,
       CODE_FROM_RAM_24,
       CODE_FROM_RAM_32,
       CODE_FROM_RAM_31,
       CODE_FROM_RAM_28,
       CODE_FROM_RAM_26,
       CODE_FROM_RAM_14,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_9,
       CODE_FROM_RAM_7,
       CODE_FROM_RAM_16,
       CODE_FROM_RAM_35,
       CODE_FROM_RAM_19
    );
output [5:5] synd_w_5;
output [3:3] synd_w;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_5;
input  CODE_FROM_RAM_21;
input  CODE_FROM_RAM_24;
input  CODE_FROM_RAM_32;
input  CODE_FROM_RAM_31;
input  CODE_FROM_RAM_28;
input  CODE_FROM_RAM_26;
input  CODE_FROM_RAM_14;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_9;
input  CODE_FROM_RAM_7;
input  CODE_FROM_RAM_16;
input  CODE_FROM_RAM_35;
input  CODE_FROM_RAM_19;

    wire \outp_0[0]_net_1 , \outp_8[0]_net_1 , \outp_2[0]_net_1 , 
        \outp_4[0]_net_1 , GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h6996) )  \outp_4[0]  (.A(\outp_2[0]_net_1 ), .B(
        CODE_FROM_RAM_16), .C(CODE_FROM_RAM_35), .D(\outp_0[0]_net_1 ), 
        .Y(\outp_4[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h6) )  \outp_0[0]  (.A(CODE_FROM_RAM_0), .B(
        CODE_FROM_RAM_5), .Y(\outp_0[0]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h6) )  \outp_5[0]  (.A(CODE_FROM_RAM_21), .B(
        CODE_FROM_RAM_24), .Y(synd_w_5[5]));
    CFG4 #( .INIT(16'h6996) )  \outp_2[0]  (.A(CODE_FROM_RAM_14), .B(
        CODE_FROM_RAM_11), .C(CODE_FROM_RAM_9), .D(CODE_FROM_RAM_7), 
        .Y(\outp_2[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(CODE_FROM_RAM_19), .B(
        \outp_4[0]_net_1 ), .C(synd_w_5[5]), .D(\outp_8[0]_net_1 ), .Y(
        synd_w[3]));
    CFG4 #( .INIT(16'h6996) )  \outp_8[0]  (.A(CODE_FROM_RAM_32), .B(
        CODE_FROM_RAM_31), .C(CODE_FROM_RAM_28), .D(CODE_FROM_RAM_26), 
        .Y(\outp_8[0]_net_1 ));
    
endmodule


module wide_xor_15s_3s_4294967295_4294967295_3s_4_2(
       synd_w_5,
       synd_w,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_5,
       CODE_FROM_RAM_21,
       CODE_FROM_RAM_24,
       CODE_FROM_RAM_32,
       CODE_FROM_RAM_31,
       CODE_FROM_RAM_28,
       CODE_FROM_RAM_26,
       CODE_FROM_RAM_14,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_9,
       CODE_FROM_RAM_7,
       CODE_FROM_RAM_16,
       CODE_FROM_RAM_35,
       CODE_FROM_RAM_19
    );
output [5:5] synd_w_5;
output [3:3] synd_w;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_5;
input  CODE_FROM_RAM_21;
input  CODE_FROM_RAM_24;
input  CODE_FROM_RAM_32;
input  CODE_FROM_RAM_31;
input  CODE_FROM_RAM_28;
input  CODE_FROM_RAM_26;
input  CODE_FROM_RAM_14;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_9;
input  CODE_FROM_RAM_7;
input  CODE_FROM_RAM_16;
input  CODE_FROM_RAM_35;
input  CODE_FROM_RAM_19;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_19 \genXOR[2].layer_xor_0  (.synd_w_5({
        synd_w_5[5]}), .synd_w({synd_w[3]}), .CODE_FROM_RAM_0(
        CODE_FROM_RAM_0), .CODE_FROM_RAM_5(CODE_FROM_RAM_5), 
        .CODE_FROM_RAM_21(CODE_FROM_RAM_21), .CODE_FROM_RAM_24(
        CODE_FROM_RAM_24), .CODE_FROM_RAM_32(CODE_FROM_RAM_32), 
        .CODE_FROM_RAM_31(CODE_FROM_RAM_31), .CODE_FROM_RAM_28(
        CODE_FROM_RAM_28), .CODE_FROM_RAM_26(CODE_FROM_RAM_26), 
        .CODE_FROM_RAM_14(CODE_FROM_RAM_14), .CODE_FROM_RAM_11(
        CODE_FROM_RAM_11), .CODE_FROM_RAM_9(CODE_FROM_RAM_9), 
        .CODE_FROM_RAM_7(CODE_FROM_RAM_7), .CODE_FROM_RAM_16(
        CODE_FROM_RAM_16), .CODE_FROM_RAM_35(CODE_FROM_RAM_35), 
        .CODE_FROM_RAM_19(CODE_FROM_RAM_19));
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_22(
       outp_9,
       outp_10,
       synd_w,
       CODE_FROM_RAM_29,
       CODE_FROM_RAM_26,
       CODE_FROM_RAM_23,
       CODE_FROM_RAM_19,
       CODE_FROM_RAM_30,
       CODE_FROM_RAM_10,
       CODE_FROM_RAM_3,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_7,
       CODE_FROM_RAM_5,
       CODE_FROM_RAM_21,
       CODE_FROM_RAM_12,
       CODE_FROM_RAM_16,
       CODE_FROM_RAM_15
    );
output [0:0] outp_9;
output [0:0] outp_10;
output [6:6] synd_w;
input  CODE_FROM_RAM_29;
input  CODE_FROM_RAM_26;
input  CODE_FROM_RAM_23;
input  CODE_FROM_RAM_19;
input  CODE_FROM_RAM_30;
input  CODE_FROM_RAM_10;
input  CODE_FROM_RAM_3;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_7;
input  CODE_FROM_RAM_5;
input  CODE_FROM_RAM_21;
input  CODE_FROM_RAM_12;
input  CODE_FROM_RAM_16;
input  CODE_FROM_RAM_15;

    wire \outp_2[0]_net_1 , \outp_4[0]_net_1 , GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h6996) )  \outp_4[0]  (.A(CODE_FROM_RAM_7), .B(
        CODE_FROM_RAM_5), .C(\outp_2[0]_net_1 ), .D(CODE_FROM_RAM_21), 
        .Y(\outp_4[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_2[0]  (.A(CODE_FROM_RAM_30), .B(
        CODE_FROM_RAM_10), .C(CODE_FROM_RAM_3), .D(CODE_FROM_RAM_0), 
        .Y(\outp_2[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp_10[0]  (.A(CODE_FROM_RAM_12), .B(
        \outp_4[0]_net_1 ), .C(CODE_FROM_RAM_16), .D(CODE_FROM_RAM_15), 
        .Y(outp_10[0]));
    CFG2 #( .INIT(4'h6) )  \outp[0]  (.A(outp_10[0]), .B(outp_9[0]), 
        .Y(synd_w[6]));
    CFG4 #( .INIT(16'h6996) )  \outp_9[0]  (.A(CODE_FROM_RAM_29), .B(
        CODE_FROM_RAM_26), .C(CODE_FROM_RAM_23), .D(CODE_FROM_RAM_19), 
        .Y(outp_9[0]));
    
endmodule


module wide_xor_15s_3s_4294967295_4294967295_3s_4_5(
       outp_9,
       outp_10,
       synd_w,
       CODE_FROM_RAM_29,
       CODE_FROM_RAM_26,
       CODE_FROM_RAM_23,
       CODE_FROM_RAM_19,
       CODE_FROM_RAM_30,
       CODE_FROM_RAM_10,
       CODE_FROM_RAM_3,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_7,
       CODE_FROM_RAM_5,
       CODE_FROM_RAM_21,
       CODE_FROM_RAM_12,
       CODE_FROM_RAM_16,
       CODE_FROM_RAM_15
    );
output [0:0] outp_9;
output [0:0] outp_10;
output [6:6] synd_w;
input  CODE_FROM_RAM_29;
input  CODE_FROM_RAM_26;
input  CODE_FROM_RAM_23;
input  CODE_FROM_RAM_19;
input  CODE_FROM_RAM_30;
input  CODE_FROM_RAM_10;
input  CODE_FROM_RAM_3;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_7;
input  CODE_FROM_RAM_5;
input  CODE_FROM_RAM_21;
input  CODE_FROM_RAM_12;
input  CODE_FROM_RAM_16;
input  CODE_FROM_RAM_15;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_22 \genXOR[2].layer_xor_0  (.outp_9({
        outp_9[0]}), .outp_10({outp_10[0]}), .synd_w({synd_w[6]}), 
        .CODE_FROM_RAM_29(CODE_FROM_RAM_29), .CODE_FROM_RAM_26(
        CODE_FROM_RAM_26), .CODE_FROM_RAM_23(CODE_FROM_RAM_23), 
        .CODE_FROM_RAM_19(CODE_FROM_RAM_19), .CODE_FROM_RAM_30(
        CODE_FROM_RAM_30), .CODE_FROM_RAM_10(CODE_FROM_RAM_10), 
        .CODE_FROM_RAM_3(CODE_FROM_RAM_3), .CODE_FROM_RAM_0(
        CODE_FROM_RAM_0), .CODE_FROM_RAM_7(CODE_FROM_RAM_7), 
        .CODE_FROM_RAM_5(CODE_FROM_RAM_5), .CODE_FROM_RAM_21(
        CODE_FROM_RAM_21), .CODE_FROM_RAM_12(CODE_FROM_RAM_12), 
        .CODE_FROM_RAM_16(CODE_FROM_RAM_16), .CODE_FROM_RAM_15(
        CODE_FROM_RAM_15));
    GND GND (.Y(GND_net_1));
    
endmodule


module 
        test_4463andcpuopration_COREEDAC_1_ham_dec_vlog_32s_7_0_4294967295_4294967295_0(
        
       COREEDAC_1_DATA_OUT,
       CODE_FROM_RAM
    );
output [31:0] COREEDAC_1_DATA_OUT;
input  [38:0] CODE_FROM_RAM;

    wire \outp_9[0] , \outp_10[0] , \synd_w[4] , N_190, \synd_w[1] , 
        \synd_w[0] , N_198, N_191, N_192, \synd_w[6] , N_205, 
        \synd_w[2] , N_188, \synd_w[3] , \synd_w[5] , N_187, N_189, 
        N_186, N_199, \err_w_0_a2_0[21]_net_1 , 
        \err_w_0_a2_1[36]_net_1 , \err_w_0_a2_0[7]_net_1 , 
        \err_w_0_a2_0[25]_net_1 , \err_w_0_a2_0[32]_net_1 , 
        \err_w_0_a2_0[34]_net_1 , N_202, N_196, \err_w_1[19] , N_206, 
        N_195, N_201, N_197, N_194, N_193, \err_w_1[37] , N_204, 
        \synd_w_5[5] , GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h78F0) )  \re_code[31]  (.A(N_191), .B(N_193), .C(
        CODE_FROM_RAM[31]), .D(N_199), .Y(COREEDAC_1_DATA_OUT[24]));
    CFG3 #( .INIT(8'h6C) )  \re_code[19]  (.A(N_197), .B(
        CODE_FROM_RAM[19]), .C(\err_w_1[19] ), .Y(
        COREEDAC_1_DATA_OUT[12]));
    CFG3 #( .INIT(8'h10) )  \err_w_0_a2_0[4]  (.A(\synd_w[2] ), .B(
        \synd_w[6] ), .C(\synd_w[4] ), .Y(N_195));
    CFG4 #( .INIT(16'h6CCC) )  \re_code[26]  (.A(N_191), .B(
        CODE_FROM_RAM[26]), .C(N_190), .D(N_194), .Y(
        COREEDAC_1_DATA_OUT[19]));
    CFG4 #( .INIT(16'h78F0) )  \re_code[15]  (.A(N_206), .B(N_190), .C(
        CODE_FROM_RAM[15]), .D(\synd_w[2] ), .Y(COREEDAC_1_DATA_OUT[8])
        );
    CFG3 #( .INIT(8'h10) )  \err_w_0_a2_2[2]  (.A(\synd_w[5] ), .B(
        \synd_w[3] ), .C(\synd_w[2] ), .Y(N_194));
    CFG4 #( .INIT(16'hF078) )  \re_code[8]  (.A(N_202), .B(N_190), .C(
        CODE_FROM_RAM[8]), .D(\synd_w[2] ), .Y(COREEDAC_1_DATA_OUT[1]));
    CFG2 #( .INIT(4'h2) )  \err_w_0_a2_0[16]  (.A(\synd_w[6] ), .B(
        \synd_w[4] ), .Y(N_205));
    CFG4 #( .INIT(16'h2000) )  \err_w_0_a2_0[34]  (.A(\synd_w[3] ), .B(
        \synd_w[1] ), .C(\synd_w[0] ), .D(\synd_w[5] ), .Y(
        \err_w_0_a2_0[34]_net_1 ));
    CFG4 #( .INIT(16'hF078) )  \re_code[18]  (.A(\err_w_1[37] ), .B(
        N_188), .C(CODE_FROM_RAM[18]), .D(\synd_w[4] ), .Y(
        COREEDAC_1_DATA_OUT[11]));
    CFG4 #( .INIT(16'h78F0) )  \re_code[29]  (.A(N_201), .B(N_205), .C(
        CODE_FROM_RAM[29]), .D(\synd_w[2] ), .Y(
        COREEDAC_1_DATA_OUT[22]));
    CFG2 #( .INIT(4'h2) )  \err_w_0_a2_1[6]  (.A(\synd_w[6] ), .B(
        \synd_w[2] ), .Y(N_188));
    CFG3 #( .INIT(8'h90) )  \err_w_0_a2_0[10]  (.A(\outp_9[0] ), .B(
        \outp_10[0] ), .C(\synd_w[4] ), .Y(N_190));
    CFG4 #( .INIT(16'h78F0) )  \re_code[25]  (.A(
        \err_w_0_a2_0[25]_net_1 ), .B(N_188), .C(CODE_FROM_RAM[25]), 
        .D(\synd_w[4] ), .Y(COREEDAC_1_DATA_OUT[18]));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h6C) )  \re_code[37]  (.A(N_197), .B(
        CODE_FROM_RAM[37]), .C(\err_w_1[37] ), .Y(
        COREEDAC_1_DATA_OUT[30]));
    CFG4 #( .INIT(16'h6AAA) )  \re_code[30]  (.A(CODE_FROM_RAM[30]), 
        .B(N_192), .C(N_187), .D(N_197), .Y(COREEDAC_1_DATA_OUT[23]));
    CFG4 #( .INIT(16'h6CCC) )  \re_code[33]  (.A(N_192), .B(
        CODE_FROM_RAM[33]), .C(N_190), .D(N_194), .Y(
        COREEDAC_1_DATA_OUT[26]));
    CFG2 #( .INIT(4'h2) )  \err_w_0_a2_0[1]  (.A(\synd_w[1] ), .B(
        \synd_w[0] ), .Y(N_191));
    CFG3 #( .INIT(8'h6C) )  \re_code[34]  (.A(N_193), .B(
        CODE_FROM_RAM[34]), .C(\err_w_0_a2_0[34]_net_1 ), .Y(
        COREEDAC_1_DATA_OUT[27]));
    CFG4 #( .INIT(16'h78F0) )  \re_code[28]  (.A(N_186), .B(N_195), .C(
        CODE_FROM_RAM[28]), .D(N_198), .Y(COREEDAC_1_DATA_OUT[21]));
    wide_xor_15s_3s_4294967295_4294967295_3s_4_1 wide_xor_2 (.synd_w({
        \synd_w[2] }), .CODE_FROM_RAM_27(CODE_FROM_RAM[29]), 
        .CODE_FROM_RAM_24(CODE_FROM_RAM[26]), .CODE_FROM_RAM_22(
        CODE_FROM_RAM[24]), .CODE_FROM_RAM_28(CODE_FROM_RAM[30]), 
        .CODE_FROM_RAM_35(CODE_FROM_RAM[37]), .CODE_FROM_RAM_14(
        CODE_FROM_RAM[16]), .CODE_FROM_RAM_10(CODE_FROM_RAM[12]), 
        .CODE_FROM_RAM_8(CODE_FROM_RAM[10]), .CODE_FROM_RAM_13(
        CODE_FROM_RAM[15]), .CODE_FROM_RAM_5(CODE_FROM_RAM[7]), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM[2]), .CODE_FROM_RAM_17(
        CODE_FROM_RAM[19]), .CODE_FROM_RAM_19(CODE_FROM_RAM[21]), 
        .CODE_FROM_RAM_34(CODE_FROM_RAM[36]), .CODE_FROM_RAM_31(
        CODE_FROM_RAM[33]));
    wide_xor_15s_3s_4294967295_4294967295_3s_4 wide_xor_0 (.synd_w({
        \synd_w[0] }), .CODE_FROM_RAM_34(CODE_FROM_RAM[34]), 
        .CODE_FROM_RAM_33(CODE_FROM_RAM[33]), .CODE_FROM_RAM_30(
        CODE_FROM_RAM[30]), .CODE_FROM_RAM_28(CODE_FROM_RAM[28]), 
        .CODE_FROM_RAM_38(CODE_FROM_RAM[38]), .CODE_FROM_RAM_16(
        CODE_FROM_RAM[16]), .CODE_FROM_RAM_14(CODE_FROM_RAM[14]), 
        .CODE_FROM_RAM_9(CODE_FROM_RAM[9]), .CODE_FROM_RAM_11(
        CODE_FROM_RAM[11]), .CODE_FROM_RAM_7(CODE_FROM_RAM[7]), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM[0]), .CODE_FROM_RAM_25(
        CODE_FROM_RAM[25]), .CODE_FROM_RAM_23(CODE_FROM_RAM[23]), 
        .CODE_FROM_RAM_19(CODE_FROM_RAM[19]), .CODE_FROM_RAM_20(
        CODE_FROM_RAM[20]));
    CFG3 #( .INIT(8'h6C) )  \re_code[12]  (.A(N_197), .B(
        CODE_FROM_RAM[12]), .C(N_204), .Y(COREEDAC_1_DATA_OUT[5]));
    CFG4 #( .INIT(16'h0100) )  \err_w_0_a2_0[5]  (.A(\synd_w[3] ), .B(
        \synd_w[1] ), .C(\synd_w[0] ), .D(\synd_w[5] ), .Y(N_206));
    wide_xor_15s_3s_4294967295_4294967295_3s_4_4 wide_xor_5 (.synd_w_5({
        \synd_w_5[5] }), .synd_w({\synd_w[5] }), .CODE_FROM_RAM_26(
        CODE_FROM_RAM[31]), .CODE_FROM_RAM_25(CODE_FROM_RAM[30]), 
        .CODE_FROM_RAM_18(CODE_FROM_RAM[23]), .CODE_FROM_RAM_15(
        CODE_FROM_RAM[20]), .CODE_FROM_RAM_32(CODE_FROM_RAM[37]), 
        .CODE_FROM_RAM_10(CODE_FROM_RAM[15]), .CODE_FROM_RAM_3(
        CODE_FROM_RAM[8]), .CODE_FROM_RAM_0(CODE_FROM_RAM[5]), 
        .CODE_FROM_RAM_8(CODE_FROM_RAM[13]), .CODE_FROM_RAM_6(
        CODE_FROM_RAM[11]), .CODE_FROM_RAM_13(CODE_FROM_RAM[18]), 
        .CODE_FROM_RAM_29(CODE_FROM_RAM[34]));
    CFG4 #( .INIT(16'h78F0) )  \re_code[36]  (.A(N_186), .B(
        \err_w_0_a2_1[36]_net_1 ), .C(CODE_FROM_RAM[36]), .D(
        \synd_w[2] ), .Y(COREEDAC_1_DATA_OUT[29]));
    CFG4 #( .INIT(16'h0200) )  \err_w_0_a2_0[8]  (.A(\synd_w[3] ), .B(
        \synd_w[1] ), .C(\synd_w[0] ), .D(\synd_w[5] ), .Y(N_202));
    wide_xor_15s_3s_4294967295_4294967295_3s_4_3 wide_xor_4 (.synd_w({
        \synd_w[4] }), .CODE_FROM_RAM_28(CODE_FROM_RAM[32]), 
        .CODE_FROM_RAM_24(CODE_FROM_RAM[28]), .CODE_FROM_RAM_22(
        CODE_FROM_RAM[26]), .CODE_FROM_RAM_21(CODE_FROM_RAM[25]), 
        .CODE_FROM_RAM_34(CODE_FROM_RAM[38]), .CODE_FROM_RAM_13(
        CODE_FROM_RAM[17]), .CODE_FROM_RAM_11(CODE_FROM_RAM[15]), 
        .CODE_FROM_RAM_9(CODE_FROM_RAM[13]), .CODE_FROM_RAM_6(
        CODE_FROM_RAM[10]), .CODE_FROM_RAM_4(CODE_FROM_RAM[8]), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM[4]), .CODE_FROM_RAM_16(
        CODE_FROM_RAM[20]), .CODE_FROM_RAM_18(CODE_FROM_RAM[22]), 
        .CODE_FROM_RAM_32(CODE_FROM_RAM[36]), .CODE_FROM_RAM_29(
        CODE_FROM_RAM[33]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h78F0) )  \re_code[22]  (.A(N_201), .B(N_188), .C(
        CODE_FROM_RAM[22]), .D(\synd_w[4] ), .Y(
        COREEDAC_1_DATA_OUT[15]));
    CFG4 #( .INIT(16'h0400) )  \err_w_0_a2_1[37]  (.A(\synd_w[3] ), .B(
        \synd_w[1] ), .C(\synd_w[0] ), .D(\synd_w[5] ), .Y(
        \err_w_1[37] ));
    CFG4 #( .INIT(16'h6AAA) )  \re_code[11]  (.A(CODE_FROM_RAM[11]), 
        .B(N_192), .C(N_187), .D(N_196), .Y(COREEDAC_1_DATA_OUT[4]));
    CFG4 #( .INIT(16'h6AAA) )  \re_code[35]  (.A(CODE_FROM_RAM[35]), 
        .B(N_191), .C(N_189), .D(N_196), .Y(COREEDAC_1_DATA_OUT[28]));
    CFG2 #( .INIT(4'h8) )  \err_w_0_a2_0[7]  (.A(\synd_w[1] ), .B(
        \synd_w[0] ), .Y(N_198));
    wide_xor_15s_3s_4294967295_4294967295_3s_4_0 wide_xor_1 (.synd_w({
        \synd_w[1] }), .CODE_FROM_RAM_34(CODE_FROM_RAM[35]), 
        .CODE_FROM_RAM_31(CODE_FROM_RAM[32]), .CODE_FROM_RAM_30(
        CODE_FROM_RAM[31]), .CODE_FROM_RAM_27(CODE_FROM_RAM[28]), 
        .CODE_FROM_RAM_36(CODE_FROM_RAM[37]), .CODE_FROM_RAM_16(
        CODE_FROM_RAM[17]), .CODE_FROM_RAM_13(CODE_FROM_RAM[14]), 
        .CODE_FROM_RAM_8(CODE_FROM_RAM[9]), .CODE_FROM_RAM_11(
        CODE_FROM_RAM[12]), .CODE_FROM_RAM_6(CODE_FROM_RAM[7]), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM[1]), .CODE_FROM_RAM_22(
        CODE_FROM_RAM[23]), .CODE_FROM_RAM_25(CODE_FROM_RAM[26]), 
        .CODE_FROM_RAM_20(CODE_FROM_RAM[21]), .CODE_FROM_RAM_17(
        CODE_FROM_RAM[18]));
    CFG4 #( .INIT(16'h78F0) )  \re_code[9]  (.A(N_186), .B(N_196), .C(
        CODE_FROM_RAM[9]), .D(N_198), .Y(COREEDAC_1_DATA_OUT[2]));
    CFG4 #( .INIT(16'hF078) )  \re_code[38]  (.A(\err_w_1[19] ), .B(
        N_190), .C(CODE_FROM_RAM[38]), .D(\synd_w[2] ), .Y(
        COREEDAC_1_DATA_OUT[31]));
    CFG4 #( .INIT(16'h78F0) )  \re_code[7]  (.A(N_186), .B(
        \err_w_0_a2_0[7]_net_1 ), .C(CODE_FROM_RAM[7]), .D(\synd_w[2] )
        , .Y(COREEDAC_1_DATA_OUT[0]));
    CFG4 #( .INIT(16'h0008) )  \err_w_0_a2_1[12]  (.A(\synd_w[3] ), .B(
        \synd_w[1] ), .C(\synd_w[0] ), .D(\synd_w[5] ), .Y(N_204));
    CFG3 #( .INIT(8'h04) )  \err_w_0_a2_0[6]  (.A(\synd_w[2] ), .B(
        \synd_w[6] ), .C(\synd_w[4] ), .Y(N_196));
    CFG4 #( .INIT(16'h78F0) )  \re_code[21]  (.A(N_186), .B(
        \err_w_0_a2_0[21]_net_1 ), .C(CODE_FROM_RAM[21]), .D(
        \synd_w[2] ), .Y(COREEDAC_1_DATA_OUT[14]));
    CFG4 #( .INIT(16'h0020) )  \err_w_0_a2_1[38]  (.A(\synd_w[3] ), .B(
        \synd_w[1] ), .C(\synd_w[0] ), .D(\synd_w[5] ), .Y(
        \err_w_1[19] ));
    CFG2 #( .INIT(4'h1) )  \err_w_0_a2_0[0]  (.A(\synd_w[3] ), .B(
        \synd_w[5] ), .Y(N_186));
    CFG4 #( .INIT(16'h0020) )  \err_w_0_a2_0_0[7]  (.A(\synd_w[0] ), 
        .B(\synd_w[4] ), .C(\synd_w[1] ), .D(\synd_w[6] ), .Y(
        \err_w_0_a2_0[7]_net_1 ));
    CFG4 #( .INIT(16'h0010) )  \err_w_0_a2_0[25]  (.A(\synd_w[3] ), .B(
        \synd_w[1] ), .C(\synd_w[0] ), .D(\synd_w[5] ), .Y(
        \err_w_0_a2_0[25]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \err_w_0_a2_0[12]  (.A(\synd_w[2] ), .B(
        \synd_w[6] ), .C(\synd_w[4] ), .Y(N_197));
    CFG4 #( .INIT(16'hF078) )  \re_code[17]  (.A(N_204), .B(N_190), .C(
        CODE_FROM_RAM[17]), .D(\synd_w[2] ), .Y(
        COREEDAC_1_DATA_OUT[10]));
    CFG4 #( .INIT(16'h78F0) )  \re_code[10]  (.A(N_201), .B(N_190), .C(
        CODE_FROM_RAM[10]), .D(\synd_w[2] ), .Y(COREEDAC_1_DATA_OUT[3])
        );
    CFG4 #( .INIT(16'h78F0) )  \re_code[13]  (.A(N_206), .B(N_188), .C(
        CODE_FROM_RAM[13]), .D(\synd_w[4] ), .Y(COREEDAC_1_DATA_OUT[6])
        );
    CFG4 #( .INIT(16'h6CCC) )  \re_code[14]  (.A(N_189), .B(
        CODE_FROM_RAM[14]), .C(N_193), .D(N_198), .Y(
        COREEDAC_1_DATA_OUT[7]));
    CFG4 #( .INIT(16'h1000) )  \err_w_0_a2_0[21]  (.A(\synd_w[0] ), .B(
        \synd_w[4] ), .C(\synd_w[1] ), .D(\synd_w[6] ), .Y(
        \err_w_0_a2_0[21]_net_1 ));
    CFG4 #( .INIT(16'h78F0) )  \re_code[32]  (.A(
        \err_w_0_a2_0[32]_net_1 ), .B(N_188), .C(CODE_FROM_RAM[32]), 
        .D(\synd_w[4] ), .Y(COREEDAC_1_DATA_OUT[25]));
    CFG4 #( .INIT(16'h0002) )  \err_w_0_a2_0[3]  (.A(\synd_w[3] ), .B(
        \synd_w[1] ), .C(\synd_w[0] ), .D(\synd_w[5] ), .Y(N_201));
    CFG3 #( .INIT(8'h01) )  \err_w_0_a2_2[0]  (.A(\synd_w[2] ), .B(
        \synd_w[6] ), .C(\synd_w[4] ), .Y(N_193));
    CFG2 #( .INIT(4'h4) )  \err_w_0_a2_1[0]  (.A(\synd_w[1] ), .B(
        \synd_w[0] ), .Y(N_192));
    CFG2 #( .INIT(4'h4) )  \err_w_0_a2_0[18]  (.A(\synd_w[3] ), .B(
        \synd_w[5] ), .Y(N_187));
    wide_xor_15s_3s_4294967295_4294967295_3s_4_2 wide_xor_3 (.synd_w_5({
        \synd_w_5[5] }), .synd_w({\synd_w[3] }), .CODE_FROM_RAM_0(
        CODE_FROM_RAM[3]), .CODE_FROM_RAM_5(CODE_FROM_RAM[8]), 
        .CODE_FROM_RAM_21(CODE_FROM_RAM[24]), .CODE_FROM_RAM_24(
        CODE_FROM_RAM[27]), .CODE_FROM_RAM_32(CODE_FROM_RAM[35]), 
        .CODE_FROM_RAM_31(CODE_FROM_RAM[34]), .CODE_FROM_RAM_28(
        CODE_FROM_RAM[31]), .CODE_FROM_RAM_26(CODE_FROM_RAM[29]), 
        .CODE_FROM_RAM_14(CODE_FROM_RAM[17]), .CODE_FROM_RAM_11(
        CODE_FROM_RAM[14]), .CODE_FROM_RAM_9(CODE_FROM_RAM[12]), 
        .CODE_FROM_RAM_7(CODE_FROM_RAM[10]), .CODE_FROM_RAM_16(
        CODE_FROM_RAM[19]), .CODE_FROM_RAM_35(CODE_FROM_RAM[38]), 
        .CODE_FROM_RAM_19(CODE_FROM_RAM[22]));
    CFG2 #( .INIT(4'h2) )  \err_w_0_a2_0[14]  (.A(\synd_w[3] ), .B(
        \synd_w[5] ), .Y(N_189));
    CFG4 #( .INIT(16'hF078) )  \re_code[27]  (.A(N_202), .B(N_188), .C(
        CODE_FROM_RAM[27]), .D(\synd_w[4] ), .Y(
        COREEDAC_1_DATA_OUT[20]));
    CFG4 #( .INIT(16'h6AAA) )  \re_code[20]  (.A(CODE_FROM_RAM[20]), 
        .B(N_192), .C(N_187), .D(N_195), .Y(COREEDAC_1_DATA_OUT[13]));
    CFG4 #( .INIT(16'h6AAA) )  \re_code[16]  (.A(CODE_FROM_RAM[16]), 
        .B(N_192), .C(N_194), .D(N_205), .Y(COREEDAC_1_DATA_OUT[9]));
    CFG4 #( .INIT(16'h0400) )  \err_w_0_a2_1[36]  (.A(\synd_w[0] ), .B(
        \synd_w[4] ), .C(\synd_w[1] ), .D(\synd_w[6] ), .Y(
        \err_w_0_a2_1[36]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \err_w_0_a2_0[31]  (.A(\synd_w[3] ), .B(
        \synd_w[5] ), .Y(N_199));
    wide_xor_15s_3s_4294967295_4294967295_3s_4_5 wide_xor_6 (.outp_9({
        \outp_9[0] }), .outp_10({\outp_10[0] }), .synd_w({\synd_w[6] })
        , .CODE_FROM_RAM_29(CODE_FROM_RAM[35]), .CODE_FROM_RAM_26(
        CODE_FROM_RAM[32]), .CODE_FROM_RAM_23(CODE_FROM_RAM[29]), 
        .CODE_FROM_RAM_19(CODE_FROM_RAM[25]), .CODE_FROM_RAM_30(
        CODE_FROM_RAM[36]), .CODE_FROM_RAM_10(CODE_FROM_RAM[16]), 
        .CODE_FROM_RAM_3(CODE_FROM_RAM[9]), .CODE_FROM_RAM_0(
        CODE_FROM_RAM[6]), .CODE_FROM_RAM_7(CODE_FROM_RAM[13]), 
        .CODE_FROM_RAM_5(CODE_FROM_RAM[11]), .CODE_FROM_RAM_21(
        CODE_FROM_RAM[27]), .CODE_FROM_RAM_12(CODE_FROM_RAM[18]), 
        .CODE_FROM_RAM_16(CODE_FROM_RAM[22]), .CODE_FROM_RAM_15(
        CODE_FROM_RAM[21]));
    CFG4 #( .INIT(16'h78F0) )  \re_code[23]  (.A(N_187), .B(N_193), .C(
        CODE_FROM_RAM[23]), .D(N_198), .Y(COREEDAC_1_DATA_OUT[16]));
    CFG3 #( .INIT(8'h6C) )  \re_code[24]  (.A(N_197), .B(
        CODE_FROM_RAM[24]), .C(N_202), .Y(COREEDAC_1_DATA_OUT[17]));
    CFG4 #( .INIT(16'h0004) )  \err_w_0_a2_0[32]  (.A(\synd_w[3] ), .B(
        \synd_w[1] ), .C(\synd_w[0] ), .D(\synd_w[5] ), .Y(
        \err_w_0_a2_0[32]_net_1 ));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_14(
       CODED_4,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_29,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_26,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_23,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_22,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_5,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_3,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_10,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_15,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_7,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_12
    );
input  [3:3] CODED_4;
output [5:5] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_29;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_26;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_23;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_22;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_5;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_3;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_10;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_15;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_7;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_12;

    wire \outp_5[0]_net_1 , \outp_4[0]_net_1 , \outp_8[0]_net_1 , 
        GND_net_1, VCC_net_1;
    
    CFG3 #( .INIT(8'h96) )  \outp_4[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_5), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_3), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_0), .Y(\outp_4[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_5[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_29), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_26), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_23), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_22), .Y(\outp_5[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_7), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_12), .C(\outp_8[0]_net_1 ), .D(
        \outp_4[0]_net_1 ), .Y(CODED[5]));
    CFG4 #( .INIT(16'h6996) )  \outp_8[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_10), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_15), .C(\outp_5[0]_net_1 ), .D(
        CODED_4[3]), .Y(\outp_8[0]_net_1 ));
    
endmodule


module wide_xor_14s_3s_4294967295_4294967295_3s_4_4(
       CODED_4,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_29,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_26,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_23,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_22,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_5,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_3,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_10,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_15,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_7,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_12
    );
input  [3:3] CODED_4;
output [5:5] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_29;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_26;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_23;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_22;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_5;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_3;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_10;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_15;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_7;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_12;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_14 \genXOR[2].layer_xor_0  (.CODED_4({
        CODED_4[3]}), .CODED({CODED[5]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_29(HDL_W_CPU_R_BUFF_0_MSG_TRP1_29)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_26(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_26), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_23(HDL_W_CPU_R_BUFF_0_MSG_TRP1_23)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_22(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_22), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_5(HDL_W_CPU_R_BUFF_0_MSG_TRP1_5), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_3(HDL_W_CPU_R_BUFF_0_MSG_TRP1_3), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1_0), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_10(HDL_W_CPU_R_BUFF_0_MSG_TRP1_10)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_15(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_15), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_7(HDL_W_CPU_R_BUFF_0_MSG_TRP1_7), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_12(HDL_W_CPU_R_BUFF_0_MSG_TRP1_12)
        );
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_11(
       CODED_1,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_27,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_26,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_11,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_6,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_23,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_20,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_19,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_16,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_14,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_5,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0
    );
input  [2:2] CODED_1;
output [2:2] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_27;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_26;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_11;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_6;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_23;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_20;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_19;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_16;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_14;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_5;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;

    wire \outp_8[0]_net_1 , \outp_7[0]_net_1 , \outp_6[0]_net_1 , 
        GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h6996) )  \outp_6[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_14), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_2), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_5), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_0), .Y(\outp_6[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_7[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_23), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_20), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_19), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_16), .Y(\outp_7[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(\outp_7[0]_net_1 ), .B(
        \outp_6[0]_net_1 ), .C(CODED_1[2]), .D(\outp_8[0]_net_1 ), .Y(
        CODED[2]));
    CFG4 #( .INIT(16'h6996) )  \outp_8[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_27), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_26), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_11), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_6), .Y(\outp_8[0]_net_1 ));
    
endmodule


module wide_xor_14s_3s_4294967295_4294967295_3s_4_1(
       CODED_1,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_27,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_26,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_11,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_6,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_23,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_20,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_19,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_16,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_14,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_5,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0
    );
input  [2:2] CODED_1;
output [2:2] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_27;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_26;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_11;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_6;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_23;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_20;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_19;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_16;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_14;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_5;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_11 \genXOR[2].layer_xor_0  (.CODED_1({
        CODED_1[2]}), .CODED({CODED[2]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_27(HDL_W_CPU_R_BUFF_0_MSG_TRP1_27)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_26(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_26), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_11(HDL_W_CPU_R_BUFF_0_MSG_TRP1_11)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_6(HDL_W_CPU_R_BUFF_0_MSG_TRP1_6)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_23(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_23), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_20(HDL_W_CPU_R_BUFF_0_MSG_TRP1_20)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_19(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_19), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_16(HDL_W_CPU_R_BUFF_0_MSG_TRP1_16)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_14(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_14), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1_2), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_5(HDL_W_CPU_R_BUFF_0_MSG_TRP1_5), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1_0));
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_10(
       CODED_2,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_16,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_14,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_11,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_24,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_10,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_25,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_28,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_30,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_19,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_21
    );
input  [3:3] CODED_2;
output [1:1] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_16;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_14;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_11;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_24;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_10;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_25;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_28;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_30;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_19;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_21;

    wire \outp_6[0]_net_1 , \outp_5[0]_net_1 , \outp_9[0]_net_1 , 
        GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h6996) )  \outp_6[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_16), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_14), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_11), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_2), .Y(\outp_6[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_5[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_24), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_10), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_0), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_25), .Y(\outp_5[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_19), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_21), .C(\outp_9[0]_net_1 ), .D(
        \outp_5[0]_net_1 ), .Y(CODED[1]));
    CFG4 #( .INIT(16'h6996) )  \outp_9[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_28), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_30), .C(\outp_6[0]_net_1 ), .D(
        CODED_2[3]), .Y(\outp_9[0]_net_1 ));
    
endmodule


module wide_xor_14s_3s_4294967295_4294967295_3s_4_0(
       CODED_2,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_16,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_14,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_11,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_24,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_10,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_25,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_28,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_30,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_19,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_21
    );
input  [3:3] CODED_2;
output [1:1] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_16;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_14;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_11;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_24;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_10;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_25;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_28;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_30;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_19;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_21;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_10 \genXOR[2].layer_xor_0  (.CODED_2({
        CODED_2[3]}), .CODED({CODED[1]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_16(HDL_W_CPU_R_BUFF_0_MSG_TRP1_16)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_14(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_14), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_11(HDL_W_CPU_R_BUFF_0_MSG_TRP1_11)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1_2)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_24(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_24), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_10(HDL_W_CPU_R_BUFF_0_MSG_TRP1_10)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1_0)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_25(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_25), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_28(HDL_W_CPU_R_BUFF_0_MSG_TRP1_28)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_30(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_30), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_19(HDL_W_CPU_R_BUFF_0_MSG_TRP1_19)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_21(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_21));
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_13(
       CODED_4,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_20,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_18,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_12,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_7,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_30,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_28,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_5,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_24,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_25,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_9
    );
input  [6:6] CODED_4;
output [4:4] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_20;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_18;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_12;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_7;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_30;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_28;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_5;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_24;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_25;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_9;

    wire \outp_5[0]_net_1 , \outp_3[0]_net_1 , \outp_7[0]_net_1 , 
        GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_3[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_30), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_28), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_5), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_0), .Y(\outp_3[0]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_7[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_24), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_25), .C(\outp_5[0]_net_1 ), .D(
        CODED_4[6]), .Y(\outp_7[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp_5[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_20), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_18), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_12), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_7), .Y(\outp_5[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_2), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_9), .C(\outp_7[0]_net_1 ), .D(
        \outp_3[0]_net_1 ), .Y(CODED[4]));
    
endmodule


module wide_xor_14s_3s_4294967295_4294967295_3s_4_3(
       CODED_4,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_20,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_18,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_12,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_7,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_30,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_28,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_5,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_24,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_25,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_9
    );
input  [6:6] CODED_4;
output [4:4] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_20;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_18;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_12;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_7;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_30;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_28;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_5;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_24;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_25;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_9;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_13 \genXOR[2].layer_xor_0  (.CODED_4({
        CODED_4[6]}), .CODED({CODED[4]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_20(HDL_W_CPU_R_BUFF_0_MSG_TRP1_20)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_18(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_18), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_12(HDL_W_CPU_R_BUFF_0_MSG_TRP1_12)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_7(HDL_W_CPU_R_BUFF_0_MSG_TRP1_7)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_30(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_30), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_28(HDL_W_CPU_R_BUFF_0_MSG_TRP1_28)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_5(HDL_W_CPU_R_BUFF_0_MSG_TRP1_5)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1_0)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_24(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_24), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_25(HDL_W_CPU_R_BUFF_0_MSG_TRP1_25)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1_2)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_9(HDL_W_CPU_R_BUFF_0_MSG_TRP1_9)
        );
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_9(
       CODED_1,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_12,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_16,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_9,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_4,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_31,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_27,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_26,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_23,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_18,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_7,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_21,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_13
    );
output [2:2] CODED_1;
output [0:0] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_12;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_16;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_9;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_4;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_31;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_27;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_26;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_23;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_18;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_7;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_21;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_13;

    wire \outp_8[0]_net_1 , \outp_7[0]_net_1 , \outp_6[0]_net_1 , 
        GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h6996) )  \outp_6[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_18), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_7), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_21), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_13), .Y(\outp_6[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_7[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_31), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_27), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_26), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_23), .Y(\outp_7[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(\outp_7[0]_net_1 ), .B(
        \outp_6[0]_net_1 ), .C(CODED_1[2]), .D(\outp_8[0]_net_1 ), .Y(
        CODED[0]));
    CFG4 #( .INIT(16'h6996) )  \outp_8[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_16), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_9), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_4), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_2), .Y(\outp_8[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \outp_1[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_0), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_12), .Y(CODED_1[2]));
    
endmodule


module wide_xor_14s_3s_4294967295_4294967295_3s_4(
       CODED_1,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_12,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_16,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_9,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_4,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_31,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_27,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_26,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_23,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_18,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_7,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_21,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_13
    );
output [2:2] CODED_1;
output [0:0] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_12;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_16;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_9;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_4;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_31;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_27;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_26;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_23;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_18;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_7;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_21;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_13;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_9 \genXOR[2].layer_xor_0  (.CODED_1({
        CODED_1[2]}), .CODED({CODED[0]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1_0), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_12(HDL_W_CPU_R_BUFF_0_MSG_TRP1_12)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_16(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_16), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_9(HDL_W_CPU_R_BUFF_0_MSG_TRP1_9), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_4(HDL_W_CPU_R_BUFF_0_MSG_TRP1_4), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1_2), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_31(HDL_W_CPU_R_BUFF_0_MSG_TRP1_31)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_27(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_27), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_26(HDL_W_CPU_R_BUFF_0_MSG_TRP1_26)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_23(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_23), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_18(HDL_W_CPU_R_BUFF_0_MSG_TRP1_18)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_7(HDL_W_CPU_R_BUFF_0_MSG_TRP1_7)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_21(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_21), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_13(HDL_W_CPU_R_BUFF_0_MSG_TRP1_13)
        );
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_15(
       CODED_4,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_13,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_16,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_23,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_20,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_12,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_9,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_7,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_4,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_26,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_18,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_27
    );
output [6:6] CODED_4;
output [6:6] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_13;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_16;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_23;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_20;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_12;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_9;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_7;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_4;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_26;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_18;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_27;

    wire \outp_7[0]_net_1 , \outp_6[0]_net_1 , \outp_5[0]_net_1 , 
        GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h6996) )  \outp_6[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_7), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_4), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_2), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_0), .Y(\outp_6[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \outp_4[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_13), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_16), .Y(CODED_4[6]));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_7[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_23), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_20), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_12), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_9), .Y(\outp_7[0]_net_1 ));
    CFG3 #( .INIT(8'h96) )  \outp_5[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_26), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_18), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_27), .Y(\outp_5[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(\outp_5[0]_net_1 ), .B(
        CODED_4[6]), .C(\outp_7[0]_net_1 ), .D(\outp_6[0]_net_1 ), .Y(
        CODED[6]));
    
endmodule


module wide_xor_14s_3s_4294967295_4294967295_3s_4_5(
       CODED_4,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_13,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_16,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_23,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_20,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_12,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_9,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_7,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_4,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_26,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_18,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_27
    );
output [6:6] CODED_4;
output [6:6] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_13;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_16;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_23;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_20;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_12;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_9;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_7;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_4;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_26;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_18;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_27;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_15 \genXOR[2].layer_xor_0  (.CODED_4({
        CODED_4[6]}), .CODED({CODED[6]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_13(HDL_W_CPU_R_BUFF_0_MSG_TRP1_13)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_16(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_16), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_23(HDL_W_CPU_R_BUFF_0_MSG_TRP1_23)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_20(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_20), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_12(HDL_W_CPU_R_BUFF_0_MSG_TRP1_12)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_9(HDL_W_CPU_R_BUFF_0_MSG_TRP1_9)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_7(HDL_W_CPU_R_BUFF_0_MSG_TRP1_7)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_4(HDL_W_CPU_R_BUFF_0_MSG_TRP1_4)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1_2)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1_0)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_26(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_26), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_18(HDL_W_CPU_R_BUFF_0_MSG_TRP1_18)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_27(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_27));
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_12(
       CODED_2,
       CODED_4,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_4,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_6,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_16,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_19,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_27,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_26,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_23,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_21,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_30,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_14,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_11,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_9,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2
    );
output [3:3] CODED_2;
output [3:3] CODED_4;
output [3:3] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_4;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_6;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_16;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_19;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_27;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_26;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_23;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_21;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_30;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_14;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_11;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_9;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;

    wire \outp_5[0]_net_1 , \outp_4[0]_net_1 , \outp_7[0]_net_1 , 
        GND_net_1, VCC_net_1;
    
    CFG2 #( .INIT(4'h6) )  \outp_4[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_16), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_19), .Y(CODED_4[3]));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_4_0[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_30), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_0), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_14), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_11), .Y(\outp_4[0]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h96) )  \outp_7[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_9), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_2), .C(\outp_4[0]_net_1 ), .Y(
        \outp_7[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \outp_5[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_27), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_26), .C(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_23), .D(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_21), .Y(\outp_5[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \outp_2[0]  (.A(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_4), .B(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_6), .Y(CODED_2[3]));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(CODED_2[3]), .B(
        CODED_4[3]), .C(\outp_7[0]_net_1 ), .D(\outp_5[0]_net_1 ), .Y(
        CODED[3]));
    
endmodule


module wide_xor_14s_3s_4294967295_4294967295_3s_4_2(
       CODED_2,
       CODED_4,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_4,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_6,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_16,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_19,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_27,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_26,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_23,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_21,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_30,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_0,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_14,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_11,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_9,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1_2
    );
output [3:3] CODED_2;
output [3:3] CODED_4;
output [3:3] CODED;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_4;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_6;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_16;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_19;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_27;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_26;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_23;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_21;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_30;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_0;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_14;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_11;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_9;
input  HDL_W_CPU_R_BUFF_0_MSG_TRP1_2;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    layer_xor_1s_3s_0_3s_1s_12 \genXOR[2].layer_xor_0  (.CODED_2({
        CODED_2[3]}), .CODED_4({CODED_4[3]}), .CODED({CODED[3]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_4(HDL_W_CPU_R_BUFF_0_MSG_TRP1_4), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_6(HDL_W_CPU_R_BUFF_0_MSG_TRP1_6), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_16(HDL_W_CPU_R_BUFF_0_MSG_TRP1_16)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_19(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_19), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_27(HDL_W_CPU_R_BUFF_0_MSG_TRP1_27)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_26(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_26), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_23(HDL_W_CPU_R_BUFF_0_MSG_TRP1_23)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_21(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_21), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_30(HDL_W_CPU_R_BUFF_0_MSG_TRP1_30)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1_0)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_14(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1_14), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_11(HDL_W_CPU_R_BUFF_0_MSG_TRP1_11)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_9(HDL_W_CPU_R_BUFF_0_MSG_TRP1_9)
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1_2)
        );
    GND GND (.Y(GND_net_1));
    
endmodule


module 
        test_4463andcpuopration_COREEDAC_1_ham_enc_vlog_32s_7_4294967295_4294967295(
        
       HDL_W_CPU_R_BUFF_0_MSG_TRP1,
       CODED
    );
input  [31:0] HDL_W_CPU_R_BUFF_0_MSG_TRP1;
output [6:0] CODED;

    wire \CODED_1[2] , \CODED_2[3] , \CODED_4[3] , \CODED_4[6] , 
        GND_net_1, VCC_net_1;
    
    wide_xor_14s_3s_4294967295_4294967295_3s_4_4 wide_xor_5 (.CODED_4({
        \CODED_4[3] }), .CODED({CODED[5]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_29(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[30]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_26(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[27]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_23(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[24]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_22(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[23]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_5(HDL_W_CPU_R_BUFF_0_MSG_TRP1[6]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_3(HDL_W_CPU_R_BUFF_0_MSG_TRP1[4]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1[1]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_10(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[11]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_15(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[16]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_7(HDL_W_CPU_R_BUFF_0_MSG_TRP1[8]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_12(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[13]));
    wide_xor_14s_3s_4294967295_4294967295_3s_4_1 wide_xor_2 (.CODED_1({
        \CODED_1[2] }), .CODED({CODED[2]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_27(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[30]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_26(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[29]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_11(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[14]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_6(HDL_W_CPU_R_BUFF_0_MSG_TRP1[9]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_23(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[26]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_20(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[23]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_19(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[22]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_16(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[19]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_14(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[17]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1[5]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_5(HDL_W_CPU_R_BUFF_0_MSG_TRP1[8]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1[3]));
    wide_xor_14s_3s_4294967295_4294967295_3s_4_0 wide_xor_1 (.CODED_2({
        \CODED_2[3] }), .CODED({CODED[1]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_16(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[16]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_14(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[14]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_11(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[11]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1[2]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_24(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[24]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_10(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[10]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1[0]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_25(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[25]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_28(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[28]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_30(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[30]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_19(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[19]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_21(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[21]));
    wide_xor_14s_3s_4294967295_4294967295_3s_4_3 wide_xor_4 (.CODED_4({
        \CODED_4[6] }), .CODED({CODED[4]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_20(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[21]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_18(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[19]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_12(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[13]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_7(HDL_W_CPU_R_BUFF_0_MSG_TRP1[8]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_30(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[31]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_28(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[29]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_5(HDL_W_CPU_R_BUFF_0_MSG_TRP1[6]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1[1]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_24(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[25]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_25(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[26]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1[3]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_9(HDL_W_CPU_R_BUFF_0_MSG_TRP1[10])
        );
    VCC VCC (.Y(VCC_net_1));
    wide_xor_14s_3s_4294967295_4294967295_3s_4 wide_xor_0 (.CODED_1({
        \CODED_1[2] }), .CODED({CODED[0]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1[0]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_12(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[12]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_16(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[16]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_9(HDL_W_CPU_R_BUFF_0_MSG_TRP1[9]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_4(HDL_W_CPU_R_BUFF_0_MSG_TRP1[4]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1[2]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_31(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[31]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_27(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[27]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_26(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[26]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_23(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[23]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_18(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[18]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_7(HDL_W_CPU_R_BUFF_0_MSG_TRP1[7]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_21(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[21]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_13(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[13]));
    GND GND (.Y(GND_net_1));
    wide_xor_14s_3s_4294967295_4294967295_3s_4_5 wide_xor_6 (.CODED_4({
        \CODED_4[6] }), .CODED({CODED[6]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_13(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[15]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_16(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[18]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_23(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[25]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_20(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[22]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_12(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[14]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_9(HDL_W_CPU_R_BUFF_0_MSG_TRP1[11])
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_7(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[9]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_4(HDL_W_CPU_R_BUFF_0_MSG_TRP1[6]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(HDL_W_CPU_R_BUFF_0_MSG_TRP1[4]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1[2]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_26(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[28]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_18(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[20]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_27(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[29]));
    wide_xor_14s_3s_4294967295_4294967295_3s_4_2 wide_xor_3 (.CODED_2({
        \CODED_2[3] }), .CODED_4({\CODED_4[3] }), .CODED({CODED[3]}), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_4(HDL_W_CPU_R_BUFF_0_MSG_TRP1[5]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_6(HDL_W_CPU_R_BUFF_0_MSG_TRP1[7]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_16(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[17]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_19(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[20]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_27(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[28]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_26(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[27]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_23(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[24]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_21(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[22]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_30(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[31]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_0(HDL_W_CPU_R_BUFF_0_MSG_TRP1[1]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_14(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[15]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_11(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[12]), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1_9(HDL_W_CPU_R_BUFF_0_MSG_TRP1[10])
        , .HDL_W_CPU_R_BUFF_0_MSG_TRP1_2(
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[3]));
    
endmodule


module test_4463andcpuopration_COREEDAC_1_ecc_Z6(
       HDL_W_CPU_R_BUFF_0_MSG_TRP1,
       CODED,
       COREEDAC_1_DATA_OUT,
       CODE_FROM_RAM
    );
input  [31:0] HDL_W_CPU_R_BUFF_0_MSG_TRP1;
output [6:0] CODED;
output [31:0] COREEDAC_1_DATA_OUT;
input  [38:0] CODE_FROM_RAM;

    wire GND_net_1, VCC_net_1;
    
    
        test_4463andcpuopration_COREEDAC_1_ham_dec_vlog_32s_7_0_4294967295_4294967295_0 
        test_4463andcpuopration_COREEDAC_1_decoder_0 (
        .COREEDAC_1_DATA_OUT({COREEDAC_1_DATA_OUT[31], 
        COREEDAC_1_DATA_OUT[30], COREEDAC_1_DATA_OUT[29], 
        COREEDAC_1_DATA_OUT[28], COREEDAC_1_DATA_OUT[27], 
        COREEDAC_1_DATA_OUT[26], COREEDAC_1_DATA_OUT[25], 
        COREEDAC_1_DATA_OUT[24], COREEDAC_1_DATA_OUT[23], 
        COREEDAC_1_DATA_OUT[22], COREEDAC_1_DATA_OUT[21], 
        COREEDAC_1_DATA_OUT[20], COREEDAC_1_DATA_OUT[19], 
        COREEDAC_1_DATA_OUT[18], COREEDAC_1_DATA_OUT[17], 
        COREEDAC_1_DATA_OUT[16], COREEDAC_1_DATA_OUT[15], 
        COREEDAC_1_DATA_OUT[14], COREEDAC_1_DATA_OUT[13], 
        COREEDAC_1_DATA_OUT[12], COREEDAC_1_DATA_OUT[11], 
        COREEDAC_1_DATA_OUT[10], COREEDAC_1_DATA_OUT[9], 
        COREEDAC_1_DATA_OUT[8], COREEDAC_1_DATA_OUT[7], 
        COREEDAC_1_DATA_OUT[6], COREEDAC_1_DATA_OUT[5], 
        COREEDAC_1_DATA_OUT[4], COREEDAC_1_DATA_OUT[3], 
        COREEDAC_1_DATA_OUT[2], COREEDAC_1_DATA_OUT[1], 
        COREEDAC_1_DATA_OUT[0]}), .CODE_FROM_RAM({CODE_FROM_RAM[38], 
        CODE_FROM_RAM[37], CODE_FROM_RAM[36], CODE_FROM_RAM[35], 
        CODE_FROM_RAM[34], CODE_FROM_RAM[33], CODE_FROM_RAM[32], 
        CODE_FROM_RAM[31], CODE_FROM_RAM[30], CODE_FROM_RAM[29], 
        CODE_FROM_RAM[28], CODE_FROM_RAM[27], CODE_FROM_RAM[26], 
        CODE_FROM_RAM[25], CODE_FROM_RAM[24], CODE_FROM_RAM[23], 
        CODE_FROM_RAM[22], CODE_FROM_RAM[21], CODE_FROM_RAM[20], 
        CODE_FROM_RAM[19], CODE_FROM_RAM[18], CODE_FROM_RAM[17], 
        CODE_FROM_RAM[16], CODE_FROM_RAM[15], CODE_FROM_RAM[14], 
        CODE_FROM_RAM[13], CODE_FROM_RAM[12], CODE_FROM_RAM[11], 
        CODE_FROM_RAM[10], CODE_FROM_RAM[9], CODE_FROM_RAM[8], 
        CODE_FROM_RAM[7], CODE_FROM_RAM[6], CODE_FROM_RAM[5], 
        CODE_FROM_RAM[4], CODE_FROM_RAM[3], CODE_FROM_RAM[2], 
        CODE_FROM_RAM[1], CODE_FROM_RAM[0]}));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
        test_4463andcpuopration_COREEDAC_1_ham_enc_vlog_32s_7_4294967295_4294967295 
        test_4463andcpuopration_COREEDAC_1_encoder_0 (
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1({HDL_W_CPU_R_BUFF_0_MSG_TRP1[31], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[30], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[29], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[28], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[27], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[26], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[25], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[24], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[23], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[22], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[21], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[20], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[19], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[18], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[17], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[16], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[15], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[14], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[13], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[12], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[11], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[10], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[9], HDL_W_CPU_R_BUFF_0_MSG_TRP1[8], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[7], HDL_W_CPU_R_BUFF_0_MSG_TRP1[6], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[5], HDL_W_CPU_R_BUFF_0_MSG_TRP1[4], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[3], HDL_W_CPU_R_BUFF_0_MSG_TRP1[2], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[1], HDL_W_CPU_R_BUFF_0_MSG_TRP1[0]})
        , .CODED({CODED[6], CODED[5], CODED[4], CODED[3], CODED[2], 
        CODED[1], CODED[0]}));
    
endmodule


module test_4463andcpuopration_COREEDAC_1_sub_edac_Z7(
       HDL_W_CPU_R_BUFF_0_MSG_TRP1,
       CODED,
       COREEDAC_1_DATA_OUT,
       CODE_FROM_RAM
    );
input  [31:0] HDL_W_CPU_R_BUFF_0_MSG_TRP1;
output [6:0] CODED;
output [31:0] COREEDAC_1_DATA_OUT;
input  [38:0] CODE_FROM_RAM;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    test_4463andcpuopration_COREEDAC_1_ecc_Z6 
        test_4463andcpuopration_COREEDAC_1_ecc_0 (
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1({HDL_W_CPU_R_BUFF_0_MSG_TRP1[31], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[30], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[29], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[28], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[27], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[26], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[25], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[24], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[23], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[22], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[21], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[20], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[19], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[18], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[17], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[16], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[15], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[14], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[13], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[12], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[11], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[10], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[9], HDL_W_CPU_R_BUFF_0_MSG_TRP1[8], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[7], HDL_W_CPU_R_BUFF_0_MSG_TRP1[6], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[5], HDL_W_CPU_R_BUFF_0_MSG_TRP1[4], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[3], HDL_W_CPU_R_BUFF_0_MSG_TRP1[2], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[1], HDL_W_CPU_R_BUFF_0_MSG_TRP1[0]})
        , .CODED({CODED[6], CODED[5], CODED[4], CODED[3], CODED[2], 
        CODED[1], CODED[0]}), .COREEDAC_1_DATA_OUT({
        COREEDAC_1_DATA_OUT[31], COREEDAC_1_DATA_OUT[30], 
        COREEDAC_1_DATA_OUT[29], COREEDAC_1_DATA_OUT[28], 
        COREEDAC_1_DATA_OUT[27], COREEDAC_1_DATA_OUT[26], 
        COREEDAC_1_DATA_OUT[25], COREEDAC_1_DATA_OUT[24], 
        COREEDAC_1_DATA_OUT[23], COREEDAC_1_DATA_OUT[22], 
        COREEDAC_1_DATA_OUT[21], COREEDAC_1_DATA_OUT[20], 
        COREEDAC_1_DATA_OUT[19], COREEDAC_1_DATA_OUT[18], 
        COREEDAC_1_DATA_OUT[17], COREEDAC_1_DATA_OUT[16], 
        COREEDAC_1_DATA_OUT[15], COREEDAC_1_DATA_OUT[14], 
        COREEDAC_1_DATA_OUT[13], COREEDAC_1_DATA_OUT[12], 
        COREEDAC_1_DATA_OUT[11], COREEDAC_1_DATA_OUT[10], 
        COREEDAC_1_DATA_OUT[9], COREEDAC_1_DATA_OUT[8], 
        COREEDAC_1_DATA_OUT[7], COREEDAC_1_DATA_OUT[6], 
        COREEDAC_1_DATA_OUT[5], COREEDAC_1_DATA_OUT[4], 
        COREEDAC_1_DATA_OUT[3], COREEDAC_1_DATA_OUT[2], 
        COREEDAC_1_DATA_OUT[1], COREEDAC_1_DATA_OUT[0]}), 
        .CODE_FROM_RAM({CODE_FROM_RAM[38], CODE_FROM_RAM[37], 
        CODE_FROM_RAM[36], CODE_FROM_RAM[35], CODE_FROM_RAM[34], 
        CODE_FROM_RAM[33], CODE_FROM_RAM[32], CODE_FROM_RAM[31], 
        CODE_FROM_RAM[30], CODE_FROM_RAM[29], CODE_FROM_RAM[28], 
        CODE_FROM_RAM[27], CODE_FROM_RAM[26], CODE_FROM_RAM[25], 
        CODE_FROM_RAM[24], CODE_FROM_RAM[23], CODE_FROM_RAM[22], 
        CODE_FROM_RAM[21], CODE_FROM_RAM[20], CODE_FROM_RAM[19], 
        CODE_FROM_RAM[18], CODE_FROM_RAM[17], CODE_FROM_RAM[16], 
        CODE_FROM_RAM[15], CODE_FROM_RAM[14], CODE_FROM_RAM[13], 
        CODE_FROM_RAM[12], CODE_FROM_RAM[11], CODE_FROM_RAM[10], 
        CODE_FROM_RAM[9], CODE_FROM_RAM[8], CODE_FROM_RAM[7], 
        CODE_FROM_RAM[6], CODE_FROM_RAM[5], CODE_FROM_RAM[4], 
        CODE_FROM_RAM[3], CODE_FROM_RAM[2], CODE_FROM_RAM[1], 
        CODE_FROM_RAM[0]}));
    
endmodule


module test_4463andcpuopration_COREEDAC_1_edac_Z8(
       HDL_W_CPU_R_BUFF_0_MSG_TRP1,
       CODED,
       COREEDAC_1_DATA_OUT,
       CODE_FROM_RAM
    );
input  [31:0] HDL_W_CPU_R_BUFF_0_MSG_TRP1;
output [6:0] CODED;
output [31:0] COREEDAC_1_DATA_OUT;
input  [38:0] CODE_FROM_RAM;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    test_4463andcpuopration_COREEDAC_1_sub_edac_Z7 
        test_4463andcpuopration_COREEDAC_1_sub_edac_0 (
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1({HDL_W_CPU_R_BUFF_0_MSG_TRP1[31], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[30], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[29], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[28], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[27], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[26], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[25], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[24], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[23], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[22], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[21], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[20], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[19], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[18], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[17], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[16], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[15], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[14], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[13], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[12], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[11], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[10], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[9], HDL_W_CPU_R_BUFF_0_MSG_TRP1[8], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[7], HDL_W_CPU_R_BUFF_0_MSG_TRP1[6], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[5], HDL_W_CPU_R_BUFF_0_MSG_TRP1[4], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[3], HDL_W_CPU_R_BUFF_0_MSG_TRP1[2], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[1], HDL_W_CPU_R_BUFF_0_MSG_TRP1[0]})
        , .CODED({CODED[6], CODED[5], CODED[4], CODED[3], CODED[2], 
        CODED[1], CODED[0]}), .COREEDAC_1_DATA_OUT({
        COREEDAC_1_DATA_OUT[31], COREEDAC_1_DATA_OUT[30], 
        COREEDAC_1_DATA_OUT[29], COREEDAC_1_DATA_OUT[28], 
        COREEDAC_1_DATA_OUT[27], COREEDAC_1_DATA_OUT[26], 
        COREEDAC_1_DATA_OUT[25], COREEDAC_1_DATA_OUT[24], 
        COREEDAC_1_DATA_OUT[23], COREEDAC_1_DATA_OUT[22], 
        COREEDAC_1_DATA_OUT[21], COREEDAC_1_DATA_OUT[20], 
        COREEDAC_1_DATA_OUT[19], COREEDAC_1_DATA_OUT[18], 
        COREEDAC_1_DATA_OUT[17], COREEDAC_1_DATA_OUT[16], 
        COREEDAC_1_DATA_OUT[15], COREEDAC_1_DATA_OUT[14], 
        COREEDAC_1_DATA_OUT[13], COREEDAC_1_DATA_OUT[12], 
        COREEDAC_1_DATA_OUT[11], COREEDAC_1_DATA_OUT[10], 
        COREEDAC_1_DATA_OUT[9], COREEDAC_1_DATA_OUT[8], 
        COREEDAC_1_DATA_OUT[7], COREEDAC_1_DATA_OUT[6], 
        COREEDAC_1_DATA_OUT[5], COREEDAC_1_DATA_OUT[4], 
        COREEDAC_1_DATA_OUT[3], COREEDAC_1_DATA_OUT[2], 
        COREEDAC_1_DATA_OUT[1], COREEDAC_1_DATA_OUT[0]}), 
        .CODE_FROM_RAM({CODE_FROM_RAM[38], CODE_FROM_RAM[37], 
        CODE_FROM_RAM[36], CODE_FROM_RAM[35], CODE_FROM_RAM[34], 
        CODE_FROM_RAM[33], CODE_FROM_RAM[32], CODE_FROM_RAM[31], 
        CODE_FROM_RAM[30], CODE_FROM_RAM[29], CODE_FROM_RAM[28], 
        CODE_FROM_RAM[27], CODE_FROM_RAM[26], CODE_FROM_RAM[25], 
        CODE_FROM_RAM[24], CODE_FROM_RAM[23], CODE_FROM_RAM[22], 
        CODE_FROM_RAM[21], CODE_FROM_RAM[20], CODE_FROM_RAM[19], 
        CODE_FROM_RAM[18], CODE_FROM_RAM[17], CODE_FROM_RAM[16], 
        CODE_FROM_RAM[15], CODE_FROM_RAM[14], CODE_FROM_RAM[13], 
        CODE_FROM_RAM[12], CODE_FROM_RAM[11], CODE_FROM_RAM[10], 
        CODE_FROM_RAM[9], CODE_FROM_RAM[8], CODE_FROM_RAM[7], 
        CODE_FROM_RAM[6], CODE_FROM_RAM[5], CODE_FROM_RAM[4], 
        CODE_FROM_RAM[3], CODE_FROM_RAM[2], CODE_FROM_RAM[1], 
        CODE_FROM_RAM[0]}));
    
endmodule


module test_4463andcpuopration_COREEDAC_1_actram(
       Glue_Logic_0_USER_RA_TRP1_1,
       CODED,
       HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1,
       CODE_FROM_RAM,
       HDL_W_CPU_R_BUFF_0_MSG_TRP1,
       OSC_0_XTLOSC_O2F,
       Glue_Logic_0_USER_REN_TRP1,
       RX_GPIO1_c,
       HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1
    );
input  [3:0] Glue_Logic_0_USER_RA_TRP1_1;
input  [6:0] CODED;
input  [3:0] HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1;
output [38:0] CODE_FROM_RAM;
input  [31:0] HDL_W_CPU_R_BUFF_0_MSG_TRP1;
input  OSC_0_XTLOSC_O2F;
input  Glue_Logic_0_USER_REN_TRP1;
input  RX_GPIO1_c;
input  HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1;

    wire VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    RAM1K18 test_4463andcpuopration_COREEDAC_1_actram_R0C1 (.A_DOUT({
        nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7, nc8, nc9, nc10, nc11, 
        nc12, nc13, nc14, nc15, nc16, nc17}), .B_DOUT({nc18, nc19, 
        nc20, nc21, nc22, nc23, nc24, nc25, nc26, nc27, nc28, nc29, 
        nc30, nc31, nc32, CODE_FROM_RAM[38], CODE_FROM_RAM[37], 
        CODE_FROM_RAM[36]}), .BUSY(), .A_CLK(OSC_0_XTLOSC_O2F), 
        .A_DOUT_CLK(VCC_net_1), .A_ARST_N(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({Glue_Logic_0_USER_REN_TRP1, VCC_net_1, 
        VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_DIN({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        Glue_Logic_0_USER_RA_TRP1_1[3], Glue_Logic_0_USER_RA_TRP1_1[2], 
        Glue_Logic_0_USER_RA_TRP1_1[1], Glue_Logic_0_USER_RA_TRP1_1[0], 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({VCC_net_1, VCC_net_1}), .B_CLK(RX_GPIO1_c), 
        .B_DOUT_CLK(VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(
        VCC_net_1), .B_BLK({HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1, 
        VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(VCC_net_1), 
        .B_DOUT_SRST_N(VCC_net_1), .B_DIN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[31], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[30], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[29]}), .B_ADDR({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[3], 
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[2], 
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[1], 
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .B_WEN({VCC_net_1, 
        VCC_net_1}), .A_EN(VCC_net_1), .A_DOUT_LAT(VCC_net_1), 
        .A_WIDTH({VCC_net_1, GND_net_1, VCC_net_1}), .A_WMODE(
        GND_net_1), .B_EN(VCC_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({
        VCC_net_1, GND_net_1, VCC_net_1}), .B_WMODE(GND_net_1), 
        .SII_LOCK(GND_net_1));
    RAM1K18 test_4463andcpuopration_COREEDAC_1_actram_R0C0 (.A_DOUT({
        CODE_FROM_RAM[35], CODE_FROM_RAM[34], CODE_FROM_RAM[33], 
        CODE_FROM_RAM[32], CODE_FROM_RAM[31], CODE_FROM_RAM[30], 
        CODE_FROM_RAM[29], CODE_FROM_RAM[28], CODE_FROM_RAM[27], 
        CODE_FROM_RAM[26], CODE_FROM_RAM[25], CODE_FROM_RAM[24], 
        CODE_FROM_RAM[23], CODE_FROM_RAM[22], CODE_FROM_RAM[21], 
        CODE_FROM_RAM[20], CODE_FROM_RAM[19], CODE_FROM_RAM[18]}), 
        .B_DOUT({CODE_FROM_RAM[17], CODE_FROM_RAM[16], 
        CODE_FROM_RAM[15], CODE_FROM_RAM[14], CODE_FROM_RAM[13], 
        CODE_FROM_RAM[12], CODE_FROM_RAM[11], CODE_FROM_RAM[10], 
        CODE_FROM_RAM[9], CODE_FROM_RAM[8], CODE_FROM_RAM[7], 
        CODE_FROM_RAM[6], CODE_FROM_RAM[5], CODE_FROM_RAM[4], 
        CODE_FROM_RAM[3], CODE_FROM_RAM[2], CODE_FROM_RAM[1], 
        CODE_FROM_RAM[0]}), .BUSY(), .A_CLK(OSC_0_XTLOSC_O2F), 
        .A_DOUT_CLK(VCC_net_1), .A_ARST_N(VCC_net_1), .A_DOUT_EN(
        VCC_net_1), .A_BLK({Glue_Logic_0_USER_REN_TRP1, VCC_net_1, 
        VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(
        VCC_net_1), .A_DIN({HDL_W_CPU_R_BUFF_0_MSG_TRP1[28], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[27], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[26], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[25], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[24], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[23], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[22], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[21], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[20], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[19], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[18], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[17], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[16], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[15], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[14], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[13], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[12], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[11]}), .A_ADDR({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        Glue_Logic_0_USER_RA_TRP1_1[3], Glue_Logic_0_USER_RA_TRP1_1[2], 
        Glue_Logic_0_USER_RA_TRP1_1[1], Glue_Logic_0_USER_RA_TRP1_1[0], 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .A_WEN({VCC_net_1, VCC_net_1}), .B_CLK(RX_GPIO1_c), 
        .B_DOUT_CLK(VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(
        VCC_net_1), .B_BLK({HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1, 
        VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(VCC_net_1), 
        .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[10], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[9], HDL_W_CPU_R_BUFF_0_MSG_TRP1[8], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[7], HDL_W_CPU_R_BUFF_0_MSG_TRP1[6], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[5], HDL_W_CPU_R_BUFF_0_MSG_TRP1[4], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[3], HDL_W_CPU_R_BUFF_0_MSG_TRP1[2], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[1], HDL_W_CPU_R_BUFF_0_MSG_TRP1[0], 
        CODED[6], CODED[5], CODED[4], CODED[3], CODED[2], CODED[1], 
        CODED[0]}), .B_ADDR({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[3], 
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[2], 
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[1], 
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .B_WEN({VCC_net_1, 
        VCC_net_1}), .A_EN(VCC_net_1), .A_DOUT_LAT(VCC_net_1), 
        .A_WIDTH({VCC_net_1, GND_net_1, VCC_net_1}), .A_WMODE(
        GND_net_1), .B_EN(VCC_net_1), .B_DOUT_LAT(VCC_net_1), .B_WIDTH({
        VCC_net_1, GND_net_1, VCC_net_1}), .B_WMODE(GND_net_1), 
        .SII_LOCK(GND_net_1));
    
endmodule


module test_4463andcpuopration_COREEDAC_1_COREEDAC_Z9(
       HDL_W_CPU_R_BUFF_0_MSG_TRP1,
       COREEDAC_1_DATA_OUT,
       Glue_Logic_0_USER_RA_TRP1_1,
       HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1,
       OSC_0_XTLOSC_O2F,
       Glue_Logic_0_USER_REN_TRP1,
       RX_GPIO1_c,
       HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1
    );
input  [31:0] HDL_W_CPU_R_BUFF_0_MSG_TRP1;
output [31:0] COREEDAC_1_DATA_OUT;
input  [3:0] Glue_Logic_0_USER_RA_TRP1_1;
input  [3:0] HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1;
input  OSC_0_XTLOSC_O2F;
input  Glue_Logic_0_USER_REN_TRP1;
input  RX_GPIO1_c;
input  HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1;

    wire \CODED[0] , \CODED[1] , \CODED[2] , \CODED[3] , \CODED[4] , 
        \CODED[5] , \CODED[6] , \CODE_FROM_RAM[0] , \CODE_FROM_RAM[1] , 
        \CODE_FROM_RAM[2] , \CODE_FROM_RAM[3] , \CODE_FROM_RAM[4] , 
        \CODE_FROM_RAM[5] , \CODE_FROM_RAM[6] , \CODE_FROM_RAM[7] , 
        \CODE_FROM_RAM[8] , \CODE_FROM_RAM[9] , \CODE_FROM_RAM[10] , 
        \CODE_FROM_RAM[11] , \CODE_FROM_RAM[12] , \CODE_FROM_RAM[13] , 
        \CODE_FROM_RAM[14] , \CODE_FROM_RAM[15] , \CODE_FROM_RAM[16] , 
        \CODE_FROM_RAM[17] , \CODE_FROM_RAM[18] , \CODE_FROM_RAM[19] , 
        \CODE_FROM_RAM[20] , \CODE_FROM_RAM[21] , \CODE_FROM_RAM[22] , 
        \CODE_FROM_RAM[23] , \CODE_FROM_RAM[24] , \CODE_FROM_RAM[25] , 
        \CODE_FROM_RAM[26] , \CODE_FROM_RAM[27] , \CODE_FROM_RAM[28] , 
        \CODE_FROM_RAM[29] , \CODE_FROM_RAM[30] , \CODE_FROM_RAM[31] , 
        \CODE_FROM_RAM[32] , \CODE_FROM_RAM[33] , \CODE_FROM_RAM[34] , 
        \CODE_FROM_RAM[35] , \CODE_FROM_RAM[36] , \CODE_FROM_RAM[37] , 
        \CODE_FROM_RAM[38] , GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    test_4463andcpuopration_COREEDAC_1_edac_Z8 
        test_4463andcpuopration_COREEDAC_1_edac_0 (
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1({HDL_W_CPU_R_BUFF_0_MSG_TRP1[31], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[30], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[29], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[28], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[27], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[26], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[25], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[24], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[23], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[22], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[21], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[20], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[19], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[18], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[17], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[16], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[15], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[14], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[13], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[12], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[11], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[10], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[9], HDL_W_CPU_R_BUFF_0_MSG_TRP1[8], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[7], HDL_W_CPU_R_BUFF_0_MSG_TRP1[6], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[5], HDL_W_CPU_R_BUFF_0_MSG_TRP1[4], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[3], HDL_W_CPU_R_BUFF_0_MSG_TRP1[2], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[1], HDL_W_CPU_R_BUFF_0_MSG_TRP1[0]})
        , .CODED({\CODED[6] , \CODED[5] , \CODED[4] , \CODED[3] , 
        \CODED[2] , \CODED[1] , \CODED[0] }), .COREEDAC_1_DATA_OUT({
        COREEDAC_1_DATA_OUT[31], COREEDAC_1_DATA_OUT[30], 
        COREEDAC_1_DATA_OUT[29], COREEDAC_1_DATA_OUT[28], 
        COREEDAC_1_DATA_OUT[27], COREEDAC_1_DATA_OUT[26], 
        COREEDAC_1_DATA_OUT[25], COREEDAC_1_DATA_OUT[24], 
        COREEDAC_1_DATA_OUT[23], COREEDAC_1_DATA_OUT[22], 
        COREEDAC_1_DATA_OUT[21], COREEDAC_1_DATA_OUT[20], 
        COREEDAC_1_DATA_OUT[19], COREEDAC_1_DATA_OUT[18], 
        COREEDAC_1_DATA_OUT[17], COREEDAC_1_DATA_OUT[16], 
        COREEDAC_1_DATA_OUT[15], COREEDAC_1_DATA_OUT[14], 
        COREEDAC_1_DATA_OUT[13], COREEDAC_1_DATA_OUT[12], 
        COREEDAC_1_DATA_OUT[11], COREEDAC_1_DATA_OUT[10], 
        COREEDAC_1_DATA_OUT[9], COREEDAC_1_DATA_OUT[8], 
        COREEDAC_1_DATA_OUT[7], COREEDAC_1_DATA_OUT[6], 
        COREEDAC_1_DATA_OUT[5], COREEDAC_1_DATA_OUT[4], 
        COREEDAC_1_DATA_OUT[3], COREEDAC_1_DATA_OUT[2], 
        COREEDAC_1_DATA_OUT[1], COREEDAC_1_DATA_OUT[0]}), 
        .CODE_FROM_RAM({\CODE_FROM_RAM[38] , \CODE_FROM_RAM[37] , 
        \CODE_FROM_RAM[36] , \CODE_FROM_RAM[35] , \CODE_FROM_RAM[34] , 
        \CODE_FROM_RAM[33] , \CODE_FROM_RAM[32] , \CODE_FROM_RAM[31] , 
        \CODE_FROM_RAM[30] , \CODE_FROM_RAM[29] , \CODE_FROM_RAM[28] , 
        \CODE_FROM_RAM[27] , \CODE_FROM_RAM[26] , \CODE_FROM_RAM[25] , 
        \CODE_FROM_RAM[24] , \CODE_FROM_RAM[23] , \CODE_FROM_RAM[22] , 
        \CODE_FROM_RAM[21] , \CODE_FROM_RAM[20] , \CODE_FROM_RAM[19] , 
        \CODE_FROM_RAM[18] , \CODE_FROM_RAM[17] , \CODE_FROM_RAM[16] , 
        \CODE_FROM_RAM[15] , \CODE_FROM_RAM[14] , \CODE_FROM_RAM[13] , 
        \CODE_FROM_RAM[12] , \CODE_FROM_RAM[11] , \CODE_FROM_RAM[10] , 
        \CODE_FROM_RAM[9] , \CODE_FROM_RAM[8] , \CODE_FROM_RAM[7] , 
        \CODE_FROM_RAM[6] , \CODE_FROM_RAM[5] , \CODE_FROM_RAM[4] , 
        \CODE_FROM_RAM[3] , \CODE_FROM_RAM[2] , \CODE_FROM_RAM[1] , 
        \CODE_FROM_RAM[0] }));
    test_4463andcpuopration_COREEDAC_1_actram 
        \lsram_g4.test_4463andcpuopration_COREEDAC_1_actram_0  (
        .Glue_Logic_0_USER_RA_TRP1_1({Glue_Logic_0_USER_RA_TRP1_1[3], 
        Glue_Logic_0_USER_RA_TRP1_1[2], Glue_Logic_0_USER_RA_TRP1_1[1], 
        Glue_Logic_0_USER_RA_TRP1_1[0]}), .CODED({\CODED[6] , 
        \CODED[5] , \CODED[4] , \CODED[3] , \CODED[2] , \CODED[1] , 
        \CODED[0] }), .HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1({
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[3], 
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[2], 
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[1], 
        HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0]}), .CODE_FROM_RAM({
        \CODE_FROM_RAM[38] , \CODE_FROM_RAM[37] , \CODE_FROM_RAM[36] , 
        \CODE_FROM_RAM[35] , \CODE_FROM_RAM[34] , \CODE_FROM_RAM[33] , 
        \CODE_FROM_RAM[32] , \CODE_FROM_RAM[31] , \CODE_FROM_RAM[30] , 
        \CODE_FROM_RAM[29] , \CODE_FROM_RAM[28] , \CODE_FROM_RAM[27] , 
        \CODE_FROM_RAM[26] , \CODE_FROM_RAM[25] , \CODE_FROM_RAM[24] , 
        \CODE_FROM_RAM[23] , \CODE_FROM_RAM[22] , \CODE_FROM_RAM[21] , 
        \CODE_FROM_RAM[20] , \CODE_FROM_RAM[19] , \CODE_FROM_RAM[18] , 
        \CODE_FROM_RAM[17] , \CODE_FROM_RAM[16] , \CODE_FROM_RAM[15] , 
        \CODE_FROM_RAM[14] , \CODE_FROM_RAM[13] , \CODE_FROM_RAM[12] , 
        \CODE_FROM_RAM[11] , \CODE_FROM_RAM[10] , \CODE_FROM_RAM[9] , 
        \CODE_FROM_RAM[8] , \CODE_FROM_RAM[7] , \CODE_FROM_RAM[6] , 
        \CODE_FROM_RAM[5] , \CODE_FROM_RAM[4] , \CODE_FROM_RAM[3] , 
        \CODE_FROM_RAM[2] , \CODE_FROM_RAM[1] , \CODE_FROM_RAM[0] }), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1({HDL_W_CPU_R_BUFF_0_MSG_TRP1[31], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[30], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[29], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[28], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[27], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[26], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[25], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[24], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[23], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[22], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[21], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[20], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[19], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[18], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[17], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[16], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[15], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[14], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[13], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[12], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[11], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[10], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[9], HDL_W_CPU_R_BUFF_0_MSG_TRP1[8], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[7], HDL_W_CPU_R_BUFF_0_MSG_TRP1[6], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[5], HDL_W_CPU_R_BUFF_0_MSG_TRP1[4], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[3], HDL_W_CPU_R_BUFF_0_MSG_TRP1[2], 
        HDL_W_CPU_R_BUFF_0_MSG_TRP1[1], HDL_W_CPU_R_BUFF_0_MSG_TRP1[0]})
        , .OSC_0_XTLOSC_O2F(OSC_0_XTLOSC_O2F), 
        .Glue_Logic_0_USER_REN_TRP1(Glue_Logic_0_USER_REN_TRP1), 
        .RX_GPIO1_c(RX_GPIO1_c), .HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1(
        HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1));
    GND GND (.Y(GND_net_1));
    
endmodule


module divider(
       Bit_Count_16dec_i_1,
       P_CLK,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       TX_GPIO1_c
    );
output [3:3] Bit_Count_16dec_i_1;
output P_CLK;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  TX_GPIO1_c;

    wire Bit_Count_2dec_net_1, 
        \Bit_Count_16dec_inferred_clock_RNI1ANC[3]_net_1 , 
        \Bit_Count_16dec[3]_net_1 , Bit_Count_2dec_i_i_0, 
        \Bit_Count_16dec[0]_net_1 , \Bit_Count_16dec_i_0[0] , 
        VCC_net_1, GND_net_1, \Bit_Count_16dec[1]_net_1 , 
        \Bit_Count_16dec_RNO[1]_net_1 , \Bit_Count_16dec[2]_net_1 , 
        \Bit_Count_16dec_RNO[2]_net_1 , \un2_Bit_Count_16dec_0_0[3] ;
    
    CLKINT Bit_Count_2dec_inferred_clock_RNI1195 (.A(
        Bit_Count_2dec_net_1), .Y(P_CLK));
    CFG4 #( .INIT(16'h6CCC) )  \Bit_Count_16dec_RNO[3]  (.A(
        \Bit_Count_16dec[0]_net_1 ), .B(\Bit_Count_16dec[3]_net_1 ), 
        .C(\Bit_Count_16dec[2]_net_1 ), .D(\Bit_Count_16dec[1]_net_1 ), 
        .Y(\un2_Bit_Count_16dec_0_0[3] ));
    GND GND (.Y(GND_net_1));
    CFG1 #( .INIT(2'h1) )  \Bit_Count_16dec_RNO[0]  (.A(
        \Bit_Count_16dec[0]_net_1 ), .Y(\Bit_Count_16dec_i_0[0] ));
    CFG3 #( .INIT(8'h6A) )  \Bit_Count_16dec_RNO[2]  (.A(
        \Bit_Count_16dec[2]_net_1 ), .B(\Bit_Count_16dec[1]_net_1 ), 
        .C(\Bit_Count_16dec[0]_net_1 ), .Y(
        \Bit_Count_16dec_RNO[2]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \Bit_Count_16dec_RNO[1]  (.A(
        \Bit_Count_16dec[0]_net_1 ), .B(\Bit_Count_16dec[1]_net_1 ), 
        .Y(\Bit_Count_16dec_RNO[1]_net_1 ));
    SLE \Bit_Count_16dec[1]  (.D(\Bit_Count_16dec_RNO[1]_net_1 ), .CLK(
        TX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Bit_Count_16dec[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE Bit_Count_2dec (.D(Bit_Count_2dec_i_i_0), .CLK(TX_GPIO1_c), 
        .EN(VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(Bit_Count_2dec_net_1));
    CLKINT \Bit_Count_16dec_inferred_clock_RNI1ANC_0[3]  (.A(
        \Bit_Count_16dec_inferred_clock_RNI1ANC[3]_net_1 ), .Y(
        Bit_Count_16dec_i_1[3]));
    SLE \Bit_Count_16dec[3]  (.D(\un2_Bit_Count_16dec_0_0[3] ), .CLK(
        TX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Bit_Count_16dec[3]_net_1 ));
    SLE \Bit_Count_16dec[2]  (.D(\Bit_Count_16dec_RNO[2]_net_1 ), .CLK(
        TX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Bit_Count_16dec[2]_net_1 ));
    SLE \Bit_Count_16dec[0]  (.D(\Bit_Count_16dec_i_0[0] ), .CLK(
        TX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Bit_Count_16dec[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  Bit_Count_2dec_RNO (.A(Bit_Count_2dec_net_1)
        , .Y(Bit_Count_2dec_i_i_0));
    CFG1 #( .INIT(2'h1) )  \Bit_Count_16dec_inferred_clock_RNI1ANC[3]  
        (.A(\Bit_Count_16dec[3]_net_1 ), .Y(
        \Bit_Count_16dec_inferred_clock_RNI1ANC[3]_net_1 ));
    
endmodule


module test_4463andcpuopration_OSC_0_OSC(
       OSC_0_XTLOSC_O2F,
       XTL
    );
output OSC_0_XTLOSC_O2F;
input  XTL;

    wire N_XTLOSC_CLKINT, N_XTLOSC_CLKOUT, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    XTLOSC_FAB I_XTLOSC_FAB (.A(N_XTLOSC_CLKOUT), .CLKOUT(
        N_XTLOSC_CLKINT));
    GND GND (.Y(GND_net_1));
    XTLOSC #( .MODE(2'h3), .FREQUENCY(16.0) )  I_XTLOSC (.XTL(XTL), 
        .CLKOUT(N_XTLOSC_CLKOUT));
    CLKINT I_XTLOSC_FAB_CLKINT (.A(N_XTLOSC_CLKINT), .Y(
        OSC_0_XTLOSC_O2F));
    
endmodule


module ASM_Generato(
       stream_0,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       P_CLK,
       ASM_OUT,
       pending,
       ENASM_i_0,
       ENASM
    );
output stream_0;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  P_CLK;
output ASM_OUT;
output pending;
input  ENASM_i_0;
input  ENASM;

    wire \stream[22]_net_1 , GND_net_1, \stream_3[22]_net_1 , 
        VCC_net_1, \stream[23]_net_1 , \stream_3[23]_net_1 , 
        \stream[24]_net_1 , \stream_3[24]_net_1 , \stream[25]_net_1 , 
        \stream_3[25]_net_1 , \stream[26]_net_1 , \stream_3[26]_net_1 , 
        \stream[27]_net_1 , \stream_3[27]_net_1 , \stream[28]_net_1 , 
        \stream_3[28]_net_1 , \stream[29]_net_1 , \stream_3[29]_net_1 , 
        \stream[30]_net_1 , \stream_3[30]_net_1 , \stream[31]_net_1 , 
        \stream_3[31]_net_1 , \stream[7]_net_1 , \stream_3[7]_net_1 , 
        \stream[8]_net_1 , \stream_3[8]_net_1 , \stream[9]_net_1 , 
        \stream_3[9]_net_1 , \stream[10]_net_1 , \stream_3[10]_net_1 , 
        \stream[11]_net_1 , \stream_3[11]_net_1 , \stream[12]_net_1 , 
        \stream_3[12]_net_1 , \stream[13]_net_1 , \stream_3[13]_net_1 , 
        \stream[14]_net_1 , \stream_3[14]_net_1 , \stream[15]_net_1 , 
        \stream_3[15]_net_1 , \stream[16]_net_1 , \stream_3[16]_net_1 , 
        \stream[17]_net_1 , \stream_3[17]_net_1 , \stream[18]_net_1 , 
        \stream_3[18]_net_1 , \stream[19]_net_1 , \stream_3[19]_net_1 , 
        \stream[20]_net_1 , \stream_3[20]_net_1 , \stream[21]_net_1 , 
        \stream_3[21]_net_1 , out_3_net_1, \stream[1]_net_1 , 
        \stream_3[1]_net_1 , \stream[2]_net_1 , \stream_3[2]_net_1 , 
        \stream[3]_net_1 , \stream_3[3]_net_1 , \stream[4]_net_1 , 
        \stream_3[4]_net_1 , \stream[5]_net_1 , \stream_3[5]_net_1 , 
        \stream[6]_net_1 , \stream_3[6]_net_1 ;
    
    CFG2 #( .INIT(4'hD) )  \stream_3[25]  (.A(ENASM), .B(
        \stream[24]_net_1 ), .Y(\stream_3[25]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[14]  (.A(ENASM), .B(
        \stream[13]_net_1 ), .Y(\stream_3[14]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[10]  (.A(ENASM), .B(
        \stream[9]_net_1 ), .Y(\stream_3[10]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[2]  (.A(ENASM), .B(
        \stream[1]_net_1 ), .Y(\stream_3[2]_net_1 ));
    SLE \stream[13]  (.D(\stream_3[13]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[13]_net_1 ));
    SLE \stream[26]  (.D(\stream_3[26]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[26]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[27]  (.A(ENASM), .B(
        \stream[26]_net_1 ), .Y(\stream_3[27]_net_1 ));
    SLE \stream[16]  (.D(\stream_3[16]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[16]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[22]  (.A(ENASM), .B(
        \stream[21]_net_1 ), .Y(\stream_3[22]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[16]  (.A(ENASM), .B(
        \stream[15]_net_1 ), .Y(\stream_3[16]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[21]  (.A(ENASM), .B(
        \stream[20]_net_1 ), .Y(\stream_3[21]_net_1 ));
    SLE \stream[5]  (.D(\stream_3[5]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[5]_net_1 ));
    SLE \stream[7]  (.D(\stream_3[7]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[7]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h8) )  \stream_3[6]  (.A(ENASM), .B(
        \stream[5]_net_1 ), .Y(\stream_3[6]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[28]  (.A(ENASM), .B(
        \stream[27]_net_1 ), .Y(\stream_3[28]_net_1 ));
    SLE \stream[30]  (.D(\stream_3[30]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[30]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[29]  (.A(ENASM), .B(
        \stream[28]_net_1 ), .Y(\stream_3[29]_net_1 ));
    SLE pending_inst_1 (.D(stream_0), .CLK(P_CLK), .EN(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ALn(VCC_net_1), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(pending));
    CFG2 #( .INIT(4'hD) )  \stream_3[23]  (.A(ENASM), .B(
        \stream[22]_net_1 ), .Y(\stream_3[23]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[31]  (.A(ENASM), .B(
        \stream[30]_net_1 ), .Y(\stream_3[31]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[15]  (.A(ENASM), .B(
        \stream[14]_net_1 ), .Y(\stream_3[15]_net_1 ));
    SLE out (.D(out_3_net_1), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(ASM_OUT));
    SLE \stream[28]  (.D(\stream_3[28]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[28]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \stream[20]  (.D(\stream_3[20]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[20]_net_1 ));
    SLE \stream[8]  (.D(\stream_3[8]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[8]_net_1 ));
    SLE \stream[2]  (.D(\stream_3[2]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[2]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[17]  (.A(ENASM), .B(
        \stream[16]_net_1 ), .Y(\stream_3[17]_net_1 ));
    SLE \stream[18]  (.D(\stream_3[18]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[18]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[4]  (.A(ENASM), .B(
        \stream[3]_net_1 ), .Y(\stream_3[4]_net_1 ));
    SLE \stream[10]  (.D(\stream_3[10]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[10]_net_1 ));
    SLE \stream[6]  (.D(\stream_3[6]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[6]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[12]  (.A(ENASM), .B(
        \stream[11]_net_1 ), .Y(\stream_3[12]_net_1 ));
    SLE \stream[1]  (.D(\stream_3[1]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[1]_net_1 ));
    SLE \stream[24]  (.D(\stream_3[24]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[24]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[24]  (.A(ENASM), .B(
        \stream[23]_net_1 ), .Y(\stream_3[24]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[11]  (.A(ENASM), .B(
        \stream[10]_net_1 ), .Y(\stream_3[11]_net_1 ));
    SLE \stream[29]  (.D(\stream_3[29]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[29]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[20]  (.A(ENASM), .B(
        \stream[19]_net_1 ), .Y(\stream_3[20]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[3]  (.A(ENASM), .B(
        \stream[2]_net_1 ), .Y(\stream_3[3]_net_1 ));
    SLE \stream[14]  (.D(\stream_3[14]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[14]_net_1 ));
    SLE \stream[19]  (.D(\stream_3[19]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[19]_net_1 ));
    SLE \stream[31]  (.D(\stream_3[31]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[31]_net_1 ));
    CFG2 #( .INIT(4'h8) )  out_3 (.A(ENASM), .B(\stream[31]_net_1 ), 
        .Y(out_3_net_1));
    SLE \stream[22]  (.D(\stream_3[22]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[22]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[26]  (.A(ENASM), .B(
        \stream[25]_net_1 ), .Y(\stream_3[26]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[7]  (.A(ENASM), .B(
        \stream[6]_net_1 ), .Y(\stream_3[7]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[18]  (.A(ENASM), .B(
        \stream[17]_net_1 ), .Y(\stream_3[18]_net_1 ));
    SLE \stream[12]  (.D(\stream_3[12]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[12]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[8]  (.A(ENASM), .B(
        \stream[7]_net_1 ), .Y(\stream_3[8]_net_1 ));
    SLE \stream[25]  (.D(\stream_3[25]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[25]_net_1 ));
    SLE \stream[21]  (.D(\stream_3[21]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[21]_net_1 ));
    SLE \stream[27]  (.D(\stream_3[27]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[27]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \stream_3[19]  (.A(ENASM), .B(
        \stream[18]_net_1 ), .Y(\stream_3[19]_net_1 ));
    SLE \stream[9]  (.D(\stream_3[9]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[9]_net_1 ));
    SLE \stream[15]  (.D(\stream_3[15]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[15]_net_1 ));
    SLE \stream[11]  (.D(\stream_3[11]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[11]_net_1 ));
    SLE \stream[0]  (.D(ENASM_i_0), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(stream_0));
    CFG2 #( .INIT(4'hD) )  \stream_3[13]  (.A(ENASM), .B(
        \stream[12]_net_1 ), .Y(\stream_3[13]_net_1 ));
    SLE \stream[17]  (.D(\stream_3[17]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[17]_net_1 ));
    SLE \stream[4]  (.D(\stream_3[4]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[30]  (.A(ENASM), .B(
        \stream[29]_net_1 ), .Y(\stream_3[30]_net_1 ));
    SLE \stream[3]  (.D(\stream_3[3]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[9]  (.A(ENASM), .B(
        \stream[8]_net_1 ), .Y(\stream_3[9]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[5]  (.A(ENASM), .B(
        \stream[4]_net_1 ), .Y(\stream_3[5]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \stream_3[1]  (.A(ENASM), .B(stream_0), .Y(
        \stream_3[1]_net_1 ));
    SLE \stream[23]  (.D(\stream_3[23]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\stream[23]_net_1 ));
    
endmodule


module parallel_to_serial(
       TM_RSENC_0_CODEOUTP,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       P_CLK,
       S_OUT_0,
       TM_RSENC_0_RDY,
       P_OUT,
       En_read_buff
    );
input  [7:0] TM_RSENC_0_CODEOUTP;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  P_CLK;
output S_OUT_0;
input  TM_RSENC_0_RDY;
output P_OUT;
output En_read_buff;

    wire \Bit_Count[0]_net_1 , GND_net_1, \un1_Bit_Count_i_0[0]_net_1 , 
        VCC_net_1, \Bit_Count[1]_net_1 , \Bit_Count_RNO[1]_net_1 , 
        \Bit_Count[2]_net_1 , \Bit_Count_RNO[2]_net_1 , N_1286_i_0, 
        En_Read_Buff_3_net_1, \bit[0]_net_1 , \bit_s[0] , 
        \bit[1]_net_1 , \bit_s[1] , \bit[2]_net_1 , \bit_s[2] , 
        \bit[3]_net_1 , \bit_s[3] , \bit[4]_net_1 , \bit_s[4] , 
        \bit[5]_net_1 , \bit_s[5] , \bit[6]_net_1 , \bit_s[6] , 
        \bit[7]_net_1 , \bit_s[7] , \bit[8]_net_1 , \bit_s[8] , 
        \bit[9]_net_1 , \bit_s[9] , \bit[10]_net_1 , \bit_s[10] , 
        \bit[11]_net_1 , \bit_s[11] , \bit[12]_net_1 , \bit_s[12] , 
        \bit[13]_net_1 , \bit_s[13] , \bit[14]_net_1 , \bit_s[14] , 
        \bit[15]_net_1 , \bit_s[15]_net_1 , bit_s_365_FCO, 
        \bit_cry[0]_net_1 , \bit_cry[1]_net_1 , \bit_cry[2]_net_1 , 
        \bit_cry[3]_net_1 , \bit_cry[4]_net_1 , \bit_cry[5]_net_1 , 
        \bit_cry[6]_net_1 , \bit_cry[7]_net_1 , \bit_cry[8]_net_1 , 
        \bit_cry[9]_net_1 , \bit_cry[10]_net_1 , \bit_cry[11]_net_1 , 
        \bit_cry[12]_net_1 , \bit_cry[13]_net_1 , \bit_cry[14]_net_1 , 
        N_1286_i_1_0, N_1286_i_1_1, N_1291, N_1420, N_1423, 
        DataO_2_6_i_m3_1_2, En_Read_Buff8lto2_0_net_1, 
        En_Read_Buff_3_3_net_1, En_Read_Buff8lto10_3_net_1, 
        En_Read_Buff8lt10, En_Read_Buff8lt15;
    
    ARI1 #( .INIT(20'h48800) )  \bit_cry[12]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[12]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[11]_net_1 ), .S(\bit_s[12] ), .Y(), .FCO(
        \bit_cry[12]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  DataO_2_2_i_m3 (.A(TM_RSENC_0_CODEOUTP[2]), 
        .B(\Bit_Count[2]_net_1 ), .C(TM_RSENC_0_CODEOUTP[6]), .Y(
        N_1420));
    SLE \bit[14]  (.D(\bit_s[14] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[14]_net_1 ));
    SLE \bit[6]  (.D(\bit_s[6] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[6]_net_1 ));
    SLE \bit[11]  (.D(\bit_s[11] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[11]_net_1 ));
    SLE EnO (.D(TM_RSENC_0_RDY), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(S_OUT_0));
    CFG4 #( .INIT(16'h0213) )  DataO_RNO_1 (.A(\Bit_Count[2]_net_1 ), 
        .B(N_1291), .C(TM_RSENC_0_CODEOUTP[4]), .D(
        TM_RSENC_0_CODEOUTP[0]), .Y(N_1286_i_1_1));
    CFG2 #( .INIT(4'h7) )  \un1_Bit_Count_i_0[0]  (.A(
        \Bit_Count[0]_net_1 ), .B(TM_RSENC_0_RDY), .Y(
        \un1_Bit_Count_i_0[0]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  DataO_RNO_2 (.A(TM_RSENC_0_CODEOUTP[3]), 
        .B(TM_RSENC_0_CODEOUTP[7]), .C(DataO_2_6_i_m3_1_2), .D(
        \Bit_Count[1]_net_1 ), .Y(N_1423));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[1]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[1]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[0]_net_1 ), .S(\bit_s[1] ), .Y(), .FCO(
        \bit_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[0]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[0]_net_1 ), .D(GND_net_1), .FCI(
        bit_s_365_FCO), .S(\bit_s[0] ), .Y(), .FCO(\bit_cry[0]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[9]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[9]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[8]_net_1 ), .S(\bit_s[9] ), .Y(), .FCO(
        \bit_cry[9]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[4]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[4]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[3]_net_1 ), .S(\bit_s[4] ), .Y(), .FCO(
        \bit_cry[4]_net_1 ));
    SLE \bit[12]  (.D(\bit_s[12] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[12]_net_1 ));
    CFG4 #( .INIT(16'hFFEF) )  En_Read_Buff_3_3 (.A(\bit[12]_net_1 ), 
        .B(\bit[11]_net_1 ), .C(TM_RSENC_0_RDY), .D(\bit[14]_net_1 ), 
        .Y(En_Read_Buff_3_3_net_1));
    SLE \Bit_Count[1]  (.D(\Bit_Count_RNO[1]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[1]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  En_Read_Buff8lto10_3 (.A(\bit[9]_net_1 )
        , .B(\bit[7]_net_1 ), .C(\bit[6]_net_1 ), .D(\bit[5]_net_1 ), 
        .Y(En_Read_Buff8lto10_3_net_1));
    SLE \bit[9]  (.D(\bit_s[9] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[9]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    SLE DataO (.D(N_1286_i_0), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(P_OUT));
    CFG2 #( .INIT(4'hE) )  \Bit_Count_RNILOHL[0]  (.A(
        \Bit_Count[1]_net_1 ), .B(\Bit_Count[0]_net_1 ), .Y(N_1291));
    CFG4 #( .INIT(16'hFEEE) )  En_Read_Buff8lto4 (.A(\bit[4]_net_1 ), 
        .B(\bit[3]_net_1 ), .C(\bit[1]_net_1 ), .D(
        En_Read_Buff8lto2_0_net_1), .Y(En_Read_Buff8lt10));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[14]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[14]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[13]_net_1 ), .S(\bit_s[14] ), .Y(), .FCO(
        \bit_cry[14]_net_1 ));
    SLE \Bit_Count[2]  (.D(\Bit_Count_RNO[2]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  En_Read_Buff8lto2_0 (.A(\bit[0]_net_1 ), .B(
        \bit[2]_net_1 ), .Y(En_Read_Buff8lto2_0_net_1));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[10]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[10]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[9]_net_1 ), .S(\bit_s[10] ), .Y(), .FCO(
        \bit_cry[10]_net_1 ));
    SLE \bit[1]  (.D(\bit_s[1] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[1]_net_1 ));
    CFG4 #( .INIT(16'h04AE) )  DataO_RNO_0 (.A(\Bit_Count[0]_net_1 ), 
        .B(\Bit_Count[1]_net_1 ), .C(N_1420), .D(N_1423), .Y(
        N_1286_i_1_0));
    GND GND (.Y(GND_net_1));
    SLE \bit[5]  (.D(\bit_s[5] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[5]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[6]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[6]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[5]_net_1 ), .S(\bit_s[6] ), .Y(), .FCO(
        \bit_cry[6]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  En_Read_Buff_3 (.A(\bit[15]_net_1 ), .B(
        \bit[13]_net_1 ), .C(En_Read_Buff_3_3_net_1), .D(
        En_Read_Buff8lt15), .Y(En_Read_Buff_3_net_1));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[5]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[5]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[4]_net_1 ), .S(\bit_s[5] ), .Y(), .FCO(
        \bit_cry[5]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[2]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[2]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[1]_net_1 ), .S(\bit_s[2] ), .Y(), .FCO(
        \bit_cry[2]_net_1 ));
    CFG3 #( .INIT(8'hD7) )  \Bit_Count_RNO[1]  (.A(TM_RSENC_0_RDY), .B(
        \Bit_Count[0]_net_1 ), .C(\Bit_Count[1]_net_1 ), .Y(
        \Bit_Count_RNO[1]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[3]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[3]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[2]_net_1 ), .S(\bit_s[3] ), .Y(), .FCO(
        \bit_cry[3]_net_1 ));
    SLE \bit[15]  (.D(\bit_s[15]_net_1 ), .CLK(P_CLK), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[15]_net_1 ));
    SLE \Bit_Count[0]  (.D(\un1_Bit_Count_i_0[0]_net_1 ), .CLK(P_CLK), 
        .EN(VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[0]_net_1 ));
    SLE \bit[10]  (.D(\bit_s[10] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[10]_net_1 ));
    SLE \bit[4]  (.D(\bit_s[4] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[4]_net_1 ));
    CFG3 #( .INIT(8'h9F) )  \Bit_Count_RNO[2]  (.A(
        \Bit_Count[2]_net_1 ), .B(N_1291), .C(TM_RSENC_0_RDY), .Y(
        \Bit_Count_RNO[2]_net_1 ));
    SLE \bit[7]  (.D(\bit_s[7] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[7]_net_1 ));
    CFG4 #( .INIT(16'h444E) )  DataO_RNO (.A(TM_RSENC_0_RDY), .B(
        TM_RSENC_0_CODEOUTP[0]), .C(N_1286_i_1_0), .D(N_1286_i_1_1), 
        .Y(N_1286_i_0));
    SLE \bit[2]  (.D(\bit_s[2] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[2]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[13]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[13]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[12]_net_1 ), .S(\bit_s[13] ), .Y(), .FCO(
        \bit_cry[13]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  bit_s_365 (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), 
        .S(), .Y(), .FCO(bit_s_365_FCO));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[8]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[8]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[7]_net_1 ), .S(\bit_s[8] ), .Y(), .FCO(
        \bit_cry[8]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[7]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[7]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[6]_net_1 ), .S(\bit_s[7] ), .Y(), .FCO(
        \bit_cry[7]_net_1 ));
    SLE \bit[8]  (.D(\bit_s[8] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[8]_net_1 ));
    SLE \bit[13]  (.D(\bit_s[13] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[13]_net_1 ));
    SLE \bit[0]  (.D(\bit_s[0] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[0]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \bit_cry[11]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[11]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[10]_net_1 ), .S(\bit_s[11] ), .Y(), .FCO(
        \bit_cry[11]_net_1 ));
    SLE En_Read_Buff (.D(En_Read_Buff_3_net_1), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(En_read_buff));
    ARI1 #( .INIT(20'h48800) )  \bit_s[15]  (.A(VCC_net_1), .B(
        TM_RSENC_0_RDY), .C(\bit[15]_net_1 ), .D(GND_net_1), .FCI(
        \bit_cry[14]_net_1 ), .S(\bit_s[15]_net_1 ), .Y(), .FCO());
    CFG4 #( .INIT(16'h0F53) )  DataO_RNO_3 (.A(TM_RSENC_0_CODEOUTP[5]), 
        .B(TM_RSENC_0_CODEOUTP[1]), .C(\Bit_Count[2]_net_1 ), .D(
        \Bit_Count[1]_net_1 ), .Y(DataO_2_6_i_m3_1_2));
    CFG4 #( .INIT(16'h8000) )  En_Read_Buff8lto10 (.A(\bit[10]_net_1 ), 
        .B(\bit[8]_net_1 ), .C(En_Read_Buff8lto10_3_net_1), .D(
        En_Read_Buff8lt10), .Y(En_Read_Buff8lt15));
    SLE \bit[3]  (.D(\bit_s[3] ), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \bit[3]_net_1 ));
    
endmodule


module CLTU(
       CLTU_0_TC_Packet_Counter,
       CLTU_0_TC_Error_Counter,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       RX_GPIO1_c,
       CLTU_0_IP_END,
       A_1,
       ENASM_0,
       CLTU_0_Flag_RX_ing,
       CLTU_0_Block_ErrO,
       CCA_NIRQ_c,
       RX_GPIO0_c
    );
output [31:0] CLTU_0_TC_Packet_Counter;
output [31:0] CLTU_0_TC_Error_Counter;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  RX_GPIO1_c;
output CLTU_0_IP_END;
output A_1;
output ENASM_0;
output CLTU_0_Flag_RX_ing;
output CLTU_0_Block_ErrO;
input  CCA_NIRQ_c;
input  RX_GPIO0_c;

    wire \TC_Error_Counter_s[0] , \un6_DataO_i[0] , VCC_net_1, 
        \Start_Sequence_counter_9[0]_net_1 , GND_net_1, 
        \un6_DataO_i[1] , \Start_Sequence_counter_9[1]_net_1 , 
        \un6_DataO_i[2] , \Start_Sequence_counter_9[2]_net_1 , 
        \un6_DataO_i[3] , \Start_Sequence_counter_9[3]_net_1 , 
        \Parity_Counter[0]_net_1 , \Parity_Counter_9[0]_net_1 , 
        \Parity_Counter[1]_net_1 , \Parity_Counter_9[1]_net_1 , 
        \Parity_Counter[2]_net_1 , \Parity_Counter_9[2]_net_1 , 
        \block_counter[0]_net_1 , \block_counter_8[0]_net_1 , 
        \block_counter[1]_net_1 , \block_counter_8[1]_net_1 , 
        \block_counter[2]_net_1 , \block_counter_8[2]_net_1 , 
        \Shift_reg[43]_net_1 , N_4752_i_0, un1_DataO41_22_i_0, 
        \Shift_reg[44]_net_1 , N_4727_i_0, \Shift_reg[45]_net_1 , 
        N_4702_i_0, \Shift_reg[46]_net_1 , N_4677_i_0, 
        \Shift_reg[47]_net_1 , N_4652_i_0, \Shift_reg[48]_net_1 , 
        N_4627_i_0, \Shift_reg[49]_net_1 , N_59, \Shift_reg[50]_net_1 , 
        N_4580_i_0, \Shift_reg[51]_net_1 , N_4558_i_0, 
        \Shift_reg[52]_net_1 , N_4533_i_0, \Shift_reg[53]_net_1 , 
        N_4511_i_0, \Shift_reg[54]_net_1 , N_4489_i_0, 
        \Shift_reg[55]_net_1 , N_4464_i_0, \State2[0]_net_1 , 
        \State2_9[0] , un1_DataO41_12_i_0, \State2[1]_net_1 , 
        State2_2_sqmuxa, \Shift_reg[28]_net_1 , N_61, 
        \Shift_reg[29]_net_1 , N_4414_i_0, \Shift_reg[30]_net_1 , 
        N_4389_i_0, \Shift_reg[31]_net_1 , N_4364_i_0, 
        \Shift_reg[32]_net_1 , N_4342_i_0, \Shift_reg[33]_net_1 , 
        N_4317_i_0, \Shift_reg[34]_net_1 , N_4292_i_0, 
        \Shift_reg[35]_net_1 , N_4270_i_0, \Shift_reg[36]_net_1 , N_56, 
        \Shift_reg[37]_net_1 , N_4223_i_0, \Shift_reg[38]_net_1 , N_63, 
        \Shift_reg[39]_net_1 , N_4176_i_0, \Shift_reg[40]_net_1 , 
        N_4151_i_0, \Shift_reg[41]_net_1 , N_65, \Shift_reg[42]_net_1 , 
        N_4101_i_0, \Shift_reg[13]_net_1 , N_4079_i_0, 
        \Shift_reg[14]_net_1 , N_67, \Shift_reg[15]_net_1 , N_4032_i_0, 
        \Shift_reg[16]_net_1 , N_4007_i_0, \Shift_reg[17]_net_1 , 
        N_3982_i_0, \Shift_reg[18]_net_1 , N_3957_i_0, 
        \Shift_reg[19]_net_1 , N_3935_i_0, \Shift_reg[20]_net_1 , 
        N_3910_i_0, \Shift_reg[21]_net_1 , N_3885_i_0, 
        \Shift_reg[22]_net_1 , N_3863_i_0, \Shift_reg[23]_net_1 , 
        N_3841_i_0, \Shift_reg[24]_net_1 , N_3816_i_0, 
        \Shift_reg[25]_net_1 , N_3792_i_0, \Shift_reg[26]_net_1 , 
        N_3767_i_0, \Shift_reg[27]_net_1 , N_69, \Parity[5]_net_1 , 
        N_3720_i_0, un1_DataO41_10_i_0, \Parity[6]_net_1 , N_3700_i_0, 
        \Shift_reg[0]_net_1 , N_3677_i_0, \Shift_reg[1]_net_1 , 
        N_3652_i_0, \Shift_reg[2]_net_1 , N_3627_i_0, 
        \Shift_reg[3]_net_1 , N_3605_i_0, \Shift_reg[4]_net_1 , 
        N_3580_i_0, \Shift_reg[5]_net_1 , N_3558_i_0, 
        \Shift_reg[6]_net_1 , N_71, \Shift_reg[7]_net_1 , N_3508_i_0, 
        \Shift_reg[8]_net_1 , N_3483_i_0, \Shift_reg[9]_net_1 , N_73, 
        \Shift_reg[10]_net_1 , N_3433_i_0, \Shift_reg[11]_net_1 , 
        N_3408_i_0, \Shift_reg[12]_net_1 , N_75, 
        \Start_Buff[13]_net_1 , N_3366, un1_DataO41_26_i_0, 
        \Start_Buff[14]_net_1 , N_3356, \Start_Buff[15]_net_1 , N_3346, 
        \Syn_reg[0]_net_1 , N_3332_i_0, un1_DataO41_15_i_0, 
        \Syn_reg[1]_net_1 , N_3319_i_0, \Syn_reg[2]_net_1 , N_3301_i_0, 
        \Syn_reg[3]_net_1 , N_3287_i_0, \Syn_reg[4]_net_1 , N_3275_i_0, 
        \Syn_reg[5]_net_1 , N_3263_i_0, \Syn_reg[6]_net_1 , N_3245_i_0, 
        \Parity[0]_net_1 , N_3227_i_0, \Parity[1]_net_1 , N_3207_i_0, 
        \Parity[2]_net_1 , N_3187_i_0, \Parity[3]_net_1 , N_3167_i_0, 
        \Parity[4]_net_1 , N_3147_i_0, \Start_Buff[0]_net_1 , N_3132, 
        \Start_Buff[1]_net_1 , Start_Buff_10_3_380_a2_net_1, 
        \Start_Buff[2]_net_1 , N_3112, \Start_Buff[3]_net_1 , 
        Start_Buff_10_5_358_a2_net_1, \Start_Buff[4]_net_1 , N_3092, 
        \Start_Buff[5]_net_1 , N_3082, \Start_Buff[6]_net_1 , N_3072, 
        \Start_Buff[7]_net_1 , N_3062, \Start_Buff[8]_net_1 , N_3052, 
        \Start_Buff[9]_net_1 , N_3042, \Start_Buff[10]_net_1 , N_3032, 
        \Start_Buff[11]_net_1 , N_3022, \Start_Buff[12]_net_1 , 
        Start_Buff_10_14_259_a2_net_1, N_3002, un1_DataO41_19_i_0, 
        DataO_10, un1_DataO41_14_i_0, \Shift_Bit_Counter_cry_cy_Y[0] , 
        un1_DataO41_8_i_0, \State1[0]_net_1 , \State1_ns[0] , N_2992, 
        un1_DataO41_27_i_0, N_74, Flag_once_net_1, N_2969_i_0, N_88, 
        un14lto0, \Bit_Counter_lm[0] , un1_DataO41_5_i_0, 
        \Bit_Counter[1]_net_1 , \Bit_Counter_lm[1] , 
        \Bit_Counter[2]_net_1 , \Bit_Counter_lm[2] , 
        \Bit_Counter[3]_net_1 , \Bit_Counter_lm[3] , un14lto4, 
        \Bit_Counter_lm[4] , un14lto5, \Bit_Counter_lm[5] , 
        \TC_Packet_Counter_s[0] , N_295, \TC_Packet_Counter_s[1] , 
        \TC_Packet_Counter_s[2] , \TC_Packet_Counter_s[3] , 
        \TC_Packet_Counter_s[4] , \TC_Packet_Counter_s[5] , 
        \TC_Packet_Counter_s[6] , \TC_Packet_Counter_s[7] , 
        \TC_Packet_Counter_s[8] , \TC_Packet_Counter_s[9] , 
        \TC_Packet_Counter_s[10] , \TC_Packet_Counter_s[11] , 
        \TC_Packet_Counter_s[12] , \TC_Packet_Counter_s[13] , 
        \TC_Packet_Counter_s[14] , \TC_Packet_Counter_s[15] , 
        \TC_Packet_Counter_s[16] , \TC_Packet_Counter_s[17] , 
        \TC_Packet_Counter_s[18] , \TC_Packet_Counter_s[19] , 
        \TC_Packet_Counter_s[20] , \TC_Packet_Counter_s[21] , 
        \TC_Packet_Counter_s[22] , \TC_Packet_Counter_s[23] , 
        \TC_Packet_Counter_s[24] , \TC_Packet_Counter_s[25] , 
        \TC_Packet_Counter_s[26] , \TC_Packet_Counter_s[27] , 
        \TC_Packet_Counter_s[28] , \TC_Packet_Counter_s[29] , 
        \TC_Packet_Counter_s[30] , \TC_Packet_Counter_s[31] , N_79_i_1, 
        \TC_Error_Counter_s[1] , \TC_Error_Counter_s[2] , 
        \TC_Error_Counter_s[3] , \TC_Error_Counter_s[4] , 
        \TC_Error_Counter_s[5] , \TC_Error_Counter_s[6] , 
        \TC_Error_Counter_s[7] , \TC_Error_Counter_s[8] , 
        \TC_Error_Counter_s[9] , \TC_Error_Counter_s[10] , 
        \TC_Error_Counter_s[11] , \TC_Error_Counter_s[12] , 
        \TC_Error_Counter_s[13] , \TC_Error_Counter_s[14] , 
        \TC_Error_Counter_s[15] , \TC_Error_Counter_s[16] , 
        \TC_Error_Counter_s[17] , \TC_Error_Counter_s[18] , 
        \TC_Error_Counter_s[19] , \TC_Error_Counter_s[20] , 
        \TC_Error_Counter_s[21] , \TC_Error_Counter_s[22] , 
        \TC_Error_Counter_s[23] , \TC_Error_Counter_s[24] , 
        \TC_Error_Counter_s[25] , \TC_Error_Counter_s[26] , 
        \TC_Error_Counter_s[27] , \TC_Error_Counter_s[28] , 
        \TC_Error_Counter_s[29] , \TC_Error_Counter_s[30] , 
        \TC_Error_Counter_s[31]_net_1 , \un22_DataO_i[0] , 
        \Shift_Bit_Counter_s[0] , Shift_Bit_Countere, 
        \un22_DataO_i[1] , \Shift_Bit_Counter_s[1] , \un22_DataO_i[2] , 
        \Shift_Bit_Counter_s[2] , \Shift_Bit_Counter[3]_net_1 , 
        \Shift_Bit_Counter_s[3] , \Shift_Bit_Counter[4]_net_1 , 
        \Shift_Bit_Counter_s[4] , \Shift_Bit_Counter[5]_net_1 , 
        \Shift_Bit_Counter_s[5]_net_1 , TC_Packet_Counter_cry_cy, 
        un1_DataO41_18_1_0_RNIGFRM_Y, TC_Packet_Counter17_i_0, N_277, 
        \TC_Packet_Counter_cry[0] , \TC_Packet_Counter_cry[1] , 
        \TC_Packet_Counter_cry[2] , \TC_Packet_Counter_cry[3] , 
        \TC_Packet_Counter_cry[4] , \TC_Packet_Counter_cry[5] , 
        \TC_Packet_Counter_cry[6] , \TC_Packet_Counter_cry[7] , 
        \TC_Packet_Counter_cry[8] , \TC_Packet_Counter_cry[9] , 
        \TC_Packet_Counter_cry[10] , \TC_Packet_Counter_cry[11] , 
        \TC_Packet_Counter_cry[12] , \TC_Packet_Counter_cry[13] , 
        \TC_Packet_Counter_cry[14] , \TC_Packet_Counter_cry[15] , 
        \TC_Packet_Counter_cry[16] , \TC_Packet_Counter_cry[17] , 
        \TC_Packet_Counter_cry[18] , \TC_Packet_Counter_cry[19] , 
        \TC_Packet_Counter_cry[20] , \TC_Packet_Counter_cry[21] , 
        \TC_Packet_Counter_cry[22] , \TC_Packet_Counter_cry[23] , 
        \TC_Packet_Counter_cry[24] , \TC_Packet_Counter_cry[25] , 
        \TC_Packet_Counter_cry[26] , \TC_Packet_Counter_cry[27] , 
        \TC_Packet_Counter_cry[28] , \TC_Packet_Counter_cry[29] , 
        \TC_Packet_Counter_cry[30] , Shift_Bit_Counter_cry_cy, N_302, 
        \Shift_Bit_Counter_cry[0]_net_1 , 
        \Shift_Bit_Counter_cry[1]_net_1 , 
        \Shift_Bit_Counter_cry[2]_net_1 , 
        \Shift_Bit_Counter_cry[3]_net_1 , 
        \Shift_Bit_Counter_cry[4]_net_1 , TC_Error_Counter_s_367_FCO, 
        \TC_Error_Counter_cry[1]_net_1 , 
        \TC_Error_Counter_cry[2]_net_1 , 
        \TC_Error_Counter_cry[3]_net_1 , 
        \TC_Error_Counter_cry[4]_net_1 , 
        \TC_Error_Counter_cry[5]_net_1 , 
        \TC_Error_Counter_cry[6]_net_1 , 
        \TC_Error_Counter_cry[7]_net_1 , 
        \TC_Error_Counter_cry[8]_net_1 , 
        \TC_Error_Counter_cry[9]_net_1 , 
        \TC_Error_Counter_cry[10]_net_1 , 
        \TC_Error_Counter_cry[11]_net_1 , 
        \TC_Error_Counter_cry[12]_net_1 , 
        \TC_Error_Counter_cry[13]_net_1 , 
        \TC_Error_Counter_cry[14]_net_1 , 
        \TC_Error_Counter_cry[15]_net_1 , 
        \TC_Error_Counter_cry[16]_net_1 , 
        \TC_Error_Counter_cry[17]_net_1 , 
        \TC_Error_Counter_cry[18]_net_1 , 
        \TC_Error_Counter_cry[19]_net_1 , 
        \TC_Error_Counter_cry[20]_net_1 , 
        \TC_Error_Counter_cry[21]_net_1 , 
        \TC_Error_Counter_cry[22]_net_1 , 
        \TC_Error_Counter_cry[23]_net_1 , 
        \TC_Error_Counter_cry[24]_net_1 , 
        \TC_Error_Counter_cry[25]_net_1 , 
        \TC_Error_Counter_cry[26]_net_1 , 
        \TC_Error_Counter_cry[27]_net_1 , 
        \TC_Error_Counter_cry[28]_net_1 , 
        \TC_Error_Counter_cry[29]_net_1 , 
        \TC_Error_Counter_cry[30]_net_1 , Bit_Counter_s_369_FCO, 
        \Bit_Counter_cry[1]_net_1 , \Bit_Counter_s[1] , 
        \Bit_Counter_cry[2]_net_1 , \Bit_Counter_s[2] , 
        \Bit_Counter_cry[3]_net_1 , \Bit_Counter_s[3] , 
        \Bit_Counter_s[5]_net_1 , \Bit_Counter_cry[4]_net_1 , 
        \Bit_Counter_s[4] , N_53_i, N_1431, Shift_reg_68_sn_m72_6_am_1, 
        Shift_reg_68_sn_m59_i_x3_RNI590H_net_1, 
        \un1_Syn_reg_i_o3_0_x2_RNIDEP63[1]_net_1 , 
        Shift_reg_68_sn_N_32, Shift_reg_68_sn_N_49, Shift_reg_68_54_4, 
        N_4752_i_1, \Shift_reg_RNO_1[43]_net_1 , N_4756, 
        \Shift_reg_RNO_2[43]_net_1 , N_349_1, Shift_reg_68_sn_N_84_mux, 
        \un1_block_counter_4[0]_net_1 , Bit_Counter_3_sqmuxa, N_62, 
        Shift_reg_68_24_1637_i_0_0_N_2L1_net_1, N_82, 
        Shift_reg_68_sn_N_56, Shift_reg_68_24_1637_i_0_0_net_1, 
        N_436_1, Shift_reg_68_28_12_1_i_o2_1_net_1, N_86, 
        un1_Syn_reg_2, N_2846, N_2847, 
        un1_Syn_reg_2_0_a3_RNI6MOJ1_net_1, N_2843, 
        \State1_ns_0_o5_2[0]_net_1 , un1_TC_Packet_Counter17_3_net_1, 
        Shift_N_7_mux_2, Shift_reg_68_57_866_i_i_a2_3_1_1_net_1, N_123, 
        Shift_reg_68_57_866_i_i_a2_3_1_net_1, 
        Shift_reg_1_sqmuxa_1_i_o3_0_o2_RNIJK1N_0_net_1, 
        Shift_reg_68_1_2300_i_0_o2, N_1451_mux, N_4084, N_4079_i_1, 
        N_4080, un1_TC_Packet_Counter17_5_net_1, 
        Shift_reg_68_29_1522_i_0_net_1, N_1426_mux, N_3610, N_3605_i_1, 
        N_3606, Shift_reg_68_53_953_i_0_net_1, N_1437_mux, N_3846, 
        N_3841_i_1, N_3842, Shift_reg_68_39_1233_i_0_net_1, 
        \un1_Syn_reg[2] , \un1_Syn_reg[0] , \un1_Syn_reg[6] , N_113, 
        \Shift_reg_RNO_3[43]_net_1 , 
        Shift_reg_68_30_1493_i_i_o3_1_net_1, 
        un1_TC_Packet_Counter17_3_RNIS3QPC_net_1, N_114, Shift_m5_0, 
        Shift_reg_68_21_1723_i_i_a2_6_1_net_1, Shift_reg_68_sn_N_73, 
        N_250, Shift_reg_68_0_2328_i_a7_0_0_a3_0_a3_0_a2_1_1_net_1, 
        N_94_i, Shift_reg_68_13_1953_i_i_N_4L5_N_3L4_net_1, N_90, N_91, 
        Shift_reg_68_13_1953_i_i_N_4L5_N_4L6_net_1, 
        Shift_reg_68_13_1953_i_i_N_4L5_N_5L8_net_1, Shift_N_5, N_253, 
        Shift_reg_68_13_1953_i_i_1, un1_DataI_0_a3_a_a_a_a_a_a_0_41, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_42, 
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_x_RNO_net_1, 
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_x_net_1, Shift_m8_i_a3_0_sx_0, 
        Shift_m4_e_1_sx, Shift_m8_i_a3_0, 
        Shift_reg_68_0_2328_i_a7_0_0_a3_0_a3_0_a2_1_1_sx_net_1, 
        Shift_m3_e_0, r_m1_e_1, \un1_Syn_reg[4] , 
        un1_DataI_0_a3_a_a_a_a_a_a_0_40, 
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_sx_net_1, 
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_net_1, 
        Shift_reg_68_63_697_i_i_N_5L8_sx_net_1, Shift_m8_i_a3_0_sx, 
        Shift_reg_68_63_697_i_i_N_5L8_net_1, 
        Shift_reg_68_63_697_i_i_a2_0, 
        Shift_reg_68_63_697_i_i_a2_0_0_net_1, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_56, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_58, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_33, 
        un1_DataI_0_a3_a_a_a_a_a_a_x_net_1, 
        Shift_reg_68_sn_m72_7_ns_sx_0, N_2548, 
        Shift_reg_68_sn_m59_i_x3_RNI3Q7P3_net_1, 
        Shift_reg_68_sn_m72_6_ns_1, Shift_reg_68_sn_m72_7_ns_sx, 
        un1_Syn_reg_2_0_a3_RNINA0E1_net_1, Shift_N_7_1, 
        Shift_m3_0_sx_sx, Shift_m3_0_sx, 
        un1_DataI_0_a3_a_a_a_a_a_a_sx_net_1, un1_DataI, 
        un1_DataI_0_a3_a_a_a_a_a_a_N_3L3_net_1, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_32, 
        un1_DataI_0_a3_a_a_a_a_a_a_N_2L1_net_1, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_34, 
        un1_DataI_0_a3_a_a_a_a_a_a_N_5L7_net_1, 
        \State1_ns_0_o5_3[0]_net_1 , 
        Shift_reg_68_46_1115_i_i_N_8L17_1_net_1, N_215, 
        Shift_reg_68_46_1115_i_i_N_8L17_net_1, 
        un1_TC_Packet_Counter17_1_net_1, Shift_m3_e_3, 
        Shift_reg_68_1_2300_i_0_o2_0_RNIHMNKG_net_1, N_199_1, 
        Shift_reg_68_63_697_i_i_1_0, 
        Shift_reg_68_63_697_i_i_a2_3_0_net_1, Shift_m2_1_1, 
        Shift_m6_i_a4_1, N_2551, Shift_reg_68_13_1953_i_i_0_net_1, 
        Shift_reg_68_6_2159_i_i_a2_3_2_net_1, N_3868, N_3863_i_1_1, 
        N_3863_i_1, N_3866, N_4516, N_4511_i_1_1, N_4511_i_1, N_4514, 
        un1_Syn_reg_67_1_a6_3_0_net_1, \un1_Syn_reg[5] , N_376, 
        un1_Syn_reg_67_1_a6_2_1_net_1, 
        Shift_reg_68_26_1580_i_i_N_2L1_net_1, N_57, 
        Shift_reg_68_26_1580_i_i_N_4L6_net_1, Shift_m3_2_3, 
        Shift_reg_68_26_1580_i_i_1_1, 
        Shift_reg_68_26_1580_i_i_1_tz_net_1, 
        Shift_reg_68_13_1953_i_i_o3_0_0_net_1, 
        Shift_reg_68_26_1580_i_i_1, Shift_reg_68_35_1349_i_1_net_1, 
        N_3935_i_1, N_3940, N_1450_mux, N_346, 
        Shift_reg_68_8_2099_i_0_1_net_1, N_4558_i_1, N_1463_mux, 
        Shift_reg_68_31_1463_i_1_net_1, N_4032_i_1, N_4037, N_1472_mux, 
        Shift_reg_68_17_1839_i_1_net_1, N_4342_i_1, N_4347, N_1452_mux, 
        Shift_reg_68_56_895_i_1_net_1, N_3558_i_1, N_3563, N_1438_mux, 
        N_402, Shift_reg_68_37_1293_i_0_1_1_net_1, 
        Shift_reg_68_37_1293_i_0_1_net_1, 
        Shift_reg_68_46_1115_i_i_N_4L7_net_1, 
        Shift_reg_68_46_1115_i_i_N_7L14_net_1, 
        Shift_reg_68_46_1115_i_i_1, N_4727_i_1, N_403, 
        Shift_reg_68_1_2300_i_0_0_net_1, N_392, un1_CCA_i_0, 
        Start_Buff_0_sqmuxa_0_0_net_1, un1_DataO41_26_i_1, N_2682, 
        N_2675, DataO_6_55_i_m2_1_2, N_309, N_2659, N_2644, N_2627, 
        N_2624, DataO_2_15_1_2, DataO_2, N_2620, N_2617, N_1074, 
        DataO_6_15_1_2, N_330, N_339, N_333, N_400, DataO_6_30_1_2, 
        N_340, N_325, N_322, N_314, DataO_6_46_1_2, N_2673, N_318, 
        N_2663, DataO_6_53_am_1_1_net_1, DataO_6_53_am_net_1, 
        DataO_6_53_bm_1_1_net_1, DataO_6_53_bm_net_1, 
        DataO_6_6_i_m2_1_2, DataO_6_25_i_m3_1_2, DataO_6_44_1_2, 
        DataO_2_6_1_2, DataO_6_41_i_m2_1_2, DataO_6_10_i_m2_1_2, 
        DataO_2_10_1_2, DataO_6_18_i_m2_1_2, DataO_6_21_i_m2_1_2, 
        DataO_6_29_i_m2_0_5, DataO_6_37_i_m2_1_2, DataO_2_13_1_2, 
        DataO_2_3_1_2, DataO_6_34_1_2, DataO_6_3_i_m2_1_2, 
        DataO_6_13_i_m2_1_2, Shift_reg_68_40_1205_i_m4_am_net_1, 
        Shift_reg_68_40_1205_i_m4_bm_net_1, N_3819, 
        Shift_reg_68_33_1407_i_m4_am_net_1, 
        Shift_reg_68_33_1407_i_m4_bm_net_1, N_3985, 
        Shift_reg_68_34_1379_i_m4_am_net_1, 
        Shift_reg_68_34_1379_i_m4_bm_net_1, N_3960, 
        Shift_reg_68_16_1869_i_m4_am_net_1, 
        Shift_reg_68_16_1869_i_m4_bm_net_1, N_4367, 
        Shift_reg_68_22_1695_i_m4_am_net_1, 
        Shift_reg_68_22_1695_i_m4_bm_net_1, N_4226, 
        Shift_reg_68_25_1609_i_m4_am_net_1, 
        Shift_reg_68_25_1609_i_m4_bm_net_1, N_4154, 
        Shift_reg_68_55_925_i_m4_am_net_1, 
        Shift_reg_68_55_925_i_m4_bm_net_1, N_3583, 
        Shift_reg_68_18_1811_i_m4_am_net_1, 
        Shift_reg_68_18_1811_i_m4_bm_net_1, N_4320, 
        Shift_reg_68_51_1011_i_m4_am_net_1, 
        Shift_reg_68_51_1011_i_m4_bm_net_1, N_3655, 
        Shift_reg_68_58_838_i_m4_am_net_1, 
        Shift_reg_68_58_838_i_m4_bm_net_1, N_3511, 
        Shift_reg_68_61_754_i_m4_am_net_1, 
        Shift_reg_68_61_754_i_m4_bm_net_1, N_3436, 
        Shift_reg_68_14_1925_i_m4_am_net_1, 
        Shift_reg_68_14_1925_i_m4_bm_net_1, N_4417, 
        Shift_reg_68_27_1552_i_m4_am_net_1, 
        Shift_reg_68_27_1552_i_m4_bm_net_1, N_4104, 
        Shift_reg_68_2_2272_i_m4_am_net_1, 
        Shift_reg_68_2_2272_i_m4_bm_net_1, N_4705, 
        Shift_reg_68_3_2244_i_m4_am_net_1, 
        Shift_reg_68_3_2244_i_m4_bm_net_1, N_4680, 
        Shift_reg_68_4_2216_i_m4_am_net_1, 
        Shift_reg_68_4_2216_i_m4_bm_net_1, N_4655, 
        Shift_reg_68_59_810_i_m4_am_net_1, 
        Shift_reg_68_59_810_i_m4_bm_net_1, N_3486, 
        Shift_reg_68_52_983_i_m4_am_net_1, 
        Shift_reg_68_52_983_i_m4_bm_net_1, N_3630, 
        Shift_reg_68_42_1143_i_m4_am_net_1, 
        Shift_reg_68_42_1143_i_m4_bm_net_1, N_3770, 
        Shift_reg_68_15_1897_i_m4_am_net_1, 
        Shift_reg_68_15_1897_i_m4_bm_net_1, N_4392, 
        Shift_reg_68_62_726_i_m4_am_net_1, 
        Shift_reg_68_62_726_i_m4_bm_net_1, N_3411, 
        Shift_reg_68_32_1435_i_m4_am_net_1, 
        Shift_reg_68_32_1435_i_m4_bm_net_1, N_4010, 
        \un1_block_counter_7_am[0]_net_1 , 
        \un1_block_counter_7_bm[0]_net_1 , \un1_block_counter_7[0] , 
        Shift_reg_68_12_1982_i_m4_bm_net_1, 
        Shift_reg_68_12_1982_i_m4_am_net_1, N_4467, 
        Shift_reg_68_47_1039_i_m4_0_bm_net_1, 
        Shift_reg_68_47_1039_i_m4_0_am_net_1, N_3679, 
        \un1_Syn_reg_RNIQLBC[3]_net_1 , Shift_reg_68_sn_m47_0_ns_1, 
        \Syn_reg_RNI2RFH1[1]_net_1 , N_2176, N_118, N_206, N_4629, 
        Shift_reg_68_37_1293_i_0_o3_1_net_1, N_58, N_374, 
        Shift_reg_68_9_2070_i_0_o2_1_1_net_1, N_286, Shift_reg_68_50_2, 
        Shift_reg_68_50_5, Shift_reg_68_1_2300_i_0_o3_0_0_net_1, 
        Shift_reg_68_sn_m37_u_i_0, \Shift_reg_68_54_e_0[42] , N_1461, 
        N_101, N_1456_mux, \Shift_reg_68_54_e_1[55] , 
        Shift_m3_0_a2_2_2, Shift_reg_68_60_782_i_i_0_net_1, N_102, 
        N_210, Shift_N_7_mux_0, \State1_ns_0_a5_1_0[0]_net_1 , 
        Parity_16_1_505_i_0_o2_0_net_1, Block_ErrO_2_sqmuxa_1_i_a1_0, 
        N_21_i, un1_Start_Buff_1_5_net_1, Parity_16_3_456_i_o4_0, 
        Parity_16_5_407_i_o4_0_net_1, N_110, N_265, N_290, N_389, 
        N_356_1, Shift_reg_68_28_32_2_net_1, Shift_reg_68_28_9_2, 
        \un1_Syn_reg[3]_net_1 , Shift_reg_68_28_30_3, 
        Shift_reg_68_28_17_2, Shift_reg_68_28_29_3, N_34, N_3721, 
        N_2131_1, un1_DataO41_24_i_a3_0_1_net_1, 
        \Shift_reg_68_54_e_0[29] , \Shift_reg_68_54_e_0[7] , 
        \Shift_reg_68_54_e_0[10] , Shift_reg_68_28_28_1_net_1, 
        Shift_reg_68_28_22_1_net_1, Shift_reg_68_28_14_1, 
        Shift_reg_68_28_15_0_net_1, Shift_reg_68_28_53_0_net_1, 
        Shift_reg_68_28_11_0_net_1, Shift_reg_68_28_45_0_net_1, 
        Shift_reg_68_28_12_0_net_1, Shift_reg_68_28_51_0_net_1, 
        Shift_reg_68_28_43_0_net_1, \State1_ns_0_a5_2_6[0] , 
        \State1_ns_0_a5_2_4[0]_net_1 , un1_Start_Buff_1_6_net_1, 
        un1_Start_Buff_1_5_0, un1_Start_Buff_1_4_net_1, 
        un39_Shift_reg_0_net_1, un1_DataI_0_a3_a_a_a_a_a_a_0_46, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_45, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_44, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_43, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_38, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_37, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_36, 
        un1_DataI_0_a3_a_a_a_a_a_a_0_35, Shift_reg_68_28_25_4, 
        un1_Start_Buff_1_11_net_1, DataO_10_iv_0_a3_0_net_1, 
        Shift_reg_68_sn_N_9, N_385, N_387, N_103, N_404, N_370, 
        N_244_2, Shift_reg_68_sn_N_16, N_298, N_417_1, N_54_i, 
        Shift_reg_68_43_2, N_97_i, N_109, Shift_reg_68_sn_N_24, N_100, 
        Shift_reg_68_28_6_4, N_55, un1_block_counter_net_1, 
        \Shift_reg_68_54_e_0[4] , \Shift_reg_68_54_e_0[26] , 
        Shift_reg_68_60_782_i_i_o2_2_0_net_1, un1_DataO41_22_0_a3_0_2, 
        Shift_reg_68_28_0_0_net_1, Shift_reg_68_28_29_1_net_1, 
        Shift_reg_68_28_19_0_net_1, Shift_reg_68_28_8_0_net_1, 
        Shift_reg_68_28_9_0_net_1, Shift_reg_68_28_1_1_net_1, 
        Shift_reg_68_28_5_1_net_1, Shift_reg_68_28_32_0_net_1, 
        Shift_reg_68_28_34_0_net_1, Shift_reg_68_28_30_0_net_1, 
        Shift_reg_68_1_2300_i_0_o3_1_0_net_1, 
        Shift_reg_68_28_25_0_net_1, Shift_reg_68_28_6_0_net_1, 
        Shift_reg_68_28_17_0_net_1, Shift_reg_68_28_31_0_net_1, 
        Shift_reg_68_28_10_1_net_1, Shift_reg_68_28_35_1_net_1, 
        \State1_ns_0_a5_2_8[0]_net_1 , N_2130, N_243, 
        Shift_reg_68_sn_N_82_mux, DataO_0_sqmuxa_1_0_net_1, N_152, 
        N_398, N_357, N_2969_1, N_305, N_122, N_268, N_204, N_275, 
        N_80, N_3703, N_78, N_3190, Shift_reg_68_sn_N_50, 
        Shift_reg_68_sn_N_78_mux, N_3723, N_3150, 
        Shift_reg_68_9_2070_i_0_a3_0_0_net_1, Shift_m2_0_0, 
        un1_DataO41_24_i_a3_0_4_net_1, \Shift_reg_68_54_e_0[11] , 
        un1_DataO41_22_0_a3_0_3_net_1, \State1_ns_0_a5_2_9[0]_net_1 , 
        N_372, un1_Start_Buff_1_net_1, un1_DataO41_27_a1_0_net_1, 
        TC_Packet_Counter18_i_0, N_73_i, \Shift_reg_68_54_e_0[17] , 
        \Shift_reg_5[25]_net_1 , Shift_reg_68_sn_N_33, 
        Shift_reg_68_sn_N_42, Shift_m3_2_1, 
        Block_ErrO_0_sqmuxa_1_0_net_1, un1_State1_0_net_1, 
        Shift_reg_68_41_1171_i_a7_0, un1_State1_1_0_net_1, N_41, 
        N_3793, N_373, N_92, Shift_reg_68_50_net_1, Shift_reg_68_50_9, 
        Shift_reg_68_41_1171_i_a7_0_1_net_1, \Shift_reg_68_54_e_0[8] , 
        \Shift_reg_68_54_e_0[1] , \Shift_reg_68_54_e_0[30] , 
        Syn_reg_0_sqmuxa_0_net_1, N_354, Shift_reg_68_28_2_net_1, 
        Shift_reg_68_28_13_net_1, un1_State1_1_net_1, 
        Shift_reg_68_28_27_net_1, Shift_reg_68_28_47_net_1, 
        un1_DataO41_18_1_net_1, Shift_reg_68_28_3_4, 
        Shift_reg_68_28_42_4, N_87, Shift_reg_68_28_50_4, 
        State2_1_sqmuxa_net_1, Shift_reg_68_28_41_4, N_54, N_2188, 
        Syn_reg_0_sqmuxa_2_net_1, Start_Buff_0_sqmuxa_1_net_1, N_93, 
        N_1463, N_1466, \State1_ns_0_1[0]_net_1 , SUM_m2_1, 
        Shift_reg_68_13_1953_i_i_o3_0_0_0, un1_DataO41_22_0_0_net_1, 
        un1_DataO41_22_0_a3_1, Shift_reg_68_28_28_net_1, N_219, 
        Shift_reg_68_28_16_net_1, CO0_0, N_143, N_220, 
        Shift_reg_68_28_36_net_1, N_73_0, N_123_0, N_83, N_124, N_81, 
        N_121, N_120, N_1429_mux, N_92_0, N_85, N_105, N_75_0, N_89, 
        CO0, Shift_reg_68_41_1171_i_1_net_1, un1_DataO41_27_a0_0_net_1, 
        N_217, N_216, TC_Packet_Counter19_net_1, N_104, N_102_0, 
        un1_DataO41_1, Shift_reg_68_13_1953_i_i_1_tz_net_1, N_2121, 
        Shift_m2_0_3, Shift_reg_68_21_1723_i_i_a2_2_0_net_1, 
        Shift_reg_68_20_1753_i_a7_1_0_net_1, 
        Shift_reg_68_11_2010_i_a7_1_0_net_1, 
        Shift_reg_68_7_2129_i_a7_1_0_net_1, N_350, N_4346, N_3562, 
        N_4036, N_3939, Shift_reg_68_57_866_i_i_0_RNO_0_net_1, 
        Shift_N_9_0, N_287, Shift_reg_68_54_2, Shift_reg_68_54_net_1, 
        un1_DataO41_22_0_1_net_1, SUM_m2_e, 
        Shift_reg_68_11_2010_i_0_net_1, Shift_reg_68_7_2129_i_0_net_1, 
        Shift_reg_68_20_1753_i_0_net_1, Shift_reg_68_21_1723_i_i_a2_1, 
        Shift_reg_68_24_1637_i_0_a3_1_0_net_1, N_1445, N_1435, N_381, 
        N_272, un1_DataO41_18, Shift_reg_68_37_1293_i_0_a2_2_1_net_1, 
        Shift_reg_68_19_1783_i_0_a2_2_1_net_1, N_1433_mux, CO0_1, 
        Shift_reg_68_19_1783_i_0_0_net_1, 
        Shift_reg_68_24_1637_i_0_2_net_1, N_285, N_4494, N_4585, N_231, 
        N_171, N_4275, N_193, Shift_reg_68_57_866_i_i_0_net_1, 
        Shift_reg_68_30_1493_i_i_0_net_1, 
        Shift_reg_68_19_1783_i_0_1_net_1, 
        Shift_reg_68_37_1293_i_0_2_net_1, N_227, Shift_N_10_mux, N_172, 
        N_232, N_4630, N_3913, N_3680, N_388, 
        Shift_reg_68_11_2010_i_2_net_1, Shift_reg_68_7_2129_i_2_net_1, 
        Shift_reg_68_20_1753_i_2_net_1, Shift_reg_68_21_1723_i_i_3_1, 
        Shift_reg_68_41_1171_i_3_net_1, N_283;
    
    SLE Flag_RX_ing (.D(N_2992), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_27_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_Flag_RX_ing));
    SLE \TC_Packet_Counter[20]  (.D(\TC_Packet_Counter_s[20] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[20]));
    SLE \Shift_reg[7]  (.D(N_3508_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[7]_net_1 ));
    CFG4 #( .INIT(16'hFB40) )  Shift_reg_68_51_1011_i_m4_bm (.A(N_389), 
        .B(Shift_reg_68_28_41_4), .C(RX_GPIO0_c), .D(
        \Shift_reg[1]_net_1 ), .Y(Shift_reg_68_51_1011_i_m4_bm_net_1));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[13]  (.A(
        Shift_reg_68_28_53_0_net_1), .B(N_374), .C(RX_GPIO0_c), .D(
        \Shift_reg[13]_net_1 ), .Y(N_83));
    CFG4 #( .INIT(16'h159D) )  DataO_10_iv_0_0_RNO_27 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[7]_net_1 ), .D(\Shift_reg[3]_net_1 ), .Y(
        DataO_6_18_i_m2_1_2));
    SLE \Syn_reg[5]  (.D(N_3263_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_15_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Syn_reg[5]_net_1 ));
    CFG2 #( .INIT(4'hB) )  TC_Packet_Counter18_0_0_o2 (.A(N_277), .B(
        TC_Packet_Counter17_i_0), .Y(TC_Packet_Counter18_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[18]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[18]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[17]_net_1 ), .S(
        \TC_Error_Counter_s[18] ), .Y(), .FCO(
        \TC_Error_Counter_cry[18]_net_1 ));
    CFG4 #( .INIT(16'h0405) )  \Shift_reg_RNO[21]  (.A(
        Shift_reg_68_37_1293_i_0_1_net_1), .B(\Shift_reg[21]_net_1 ), 
        .C(Shift_reg_68_37_1293_i_0_2_net_1), .D(N_388), .Y(N_3885_i_0)
        );
    CFG4 #( .INIT(16'h2367) )  DataO_10_iv_0_0_RNO_7 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[46]_net_1 ), .D(\Shift_reg[14]_net_1 ), .Y(
        DataO_6_41_i_m2_1_2));
    CFG2 #( .INIT(4'h4) )  TC_Packet_Counter19 (.A(
        un1_TC_Packet_Counter17_1_net_1), .B(un1_DataI), .Y(
        TC_Packet_Counter19_net_1));
    CFG3 #( .INIT(8'h02) )  Shift_reg_68_63_697_i_i_1_RNO (.A(
        Shift_reg_1_sqmuxa_1_i_o3_0_o2_RNIJK1N_0_net_1), .B(
        Shift_reg_68_sn_N_56), .C(Shift_reg_68_1_2300_i_0_o2), .Y(
        Shift_m2_1_1));
    SLE \Shift_reg[3]  (.D(N_3605_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[3]_net_1 ));
    SLE \Start_Buff[1]  (.D(Start_Buff_10_3_380_a2_net_1), .CLK(
        RX_GPIO1_c), .EN(un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[1]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \Bit_Counter_lm_0[1]  (.A(
        Bit_Counter_3_sqmuxa), .B(\Bit_Counter_s[1] ), .Y(
        \Bit_Counter_lm[1] ));
    CFG3 #( .INIT(8'hA2) )  \un1_Syn_reg_i_o3_0_x2_RNITNGN[1]  (.A(
        \un1_Syn_reg[6] ), .B(N_53_i), .C(\un1_Syn_reg[0] ), .Y(
        \Shift_reg_68_54_e_0[30] ));
    CFG4 #( .INIT(16'h0F53) )  DataO_10_iv_0_a3_0_RNO_4 (.A(
        \Start_Buff[6]_net_1 ), .B(\Start_Buff[14]_net_1 ), .C(
        \un6_DataO_i[3] ), .D(\un6_DataO_i[2] ), .Y(DataO_2_10_1_2));
    CFG4 #( .INIT(16'h070F) )  Enable_RNO (.A(\State2[1]_net_1 ), .B(
        CCA_NIRQ_c), .C(un1_CCA_i_0), .D(N_305), .Y(un1_DataO41_8_i_0));
    CFG4 #( .INIT(16'h3B0A) )  Shift_reg_68_57_866_i_i_0 (.A(
        Shift_m8_i_a3_0), .B(Shift_N_5), .C(
        Shift_reg_68_57_866_i_i_0_RNO_0_net_1), .D(
        Shift_reg_68_57_866_i_i_a2_3_1_net_1), .Y(
        Shift_reg_68_57_866_i_i_0_net_1));
    CFG2 #( .INIT(4'h4) )  Shift_reg_68_28_13_2 (.A(un14lto0), .B(
        un14lto4), .Y(Shift_reg_68_28_17_2));
    CFG4 #( .INIT(16'h1007) )  Shift_reg_68_50_11 (.A(\un1_Syn_reg[2] )
        , .B(N_53_i), .C(\un1_Syn_reg[0] ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_50_2));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[42]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4104), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4101_i_0));
    CFG4 #( .INIT(16'h0400) )  Shift_reg_68_39_1233_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_93), 
        .D(N_82), .Y(N_3846));
    CFG4 #( .INIT(16'h6996) )  \Syn_reg_RNI0PFH1[0]  (.A(
        \Parity[0]_net_1 ), .B(\Syn_reg[0]_net_1 ), .C(
        \Syn_reg[6]_net_1 ), .D(\Parity[6]_net_1 ), .Y(N_1431));
    CFG2 #( .INIT(4'h8) )  Start_Buff_10_2_391_a2 (.A(N_2992), .B(
        RX_GPIO0_c), .Y(N_3132));
    CFG2 #( .INIT(4'h4) )  \un1_Start_Sequence_counter_1.CO0  (.A(
        un1_DataO41_18), .B(\un6_DataO_i[0] ), .Y(CO0_1));
    CFG4 #( .INIT(16'h32FA) )  \Shift_reg_RNO_0[22]  (.A(
        \Shift_reg[22]_net_1 ), .B(\State1[0]_net_1 ), .C(
        Shift_reg_68_sn_N_84_mux), .D(un1_TC_Packet_Counter17_5_net_1), 
        .Y(N_3863_i_1));
    CFG4 #( .INIT(16'h0F0B) )  Shift_reg_68_21_1723_i_i_a2_6_1 (.A(
        un1_TC_Packet_Counter17_3_net_1), .B(
        Shift_reg_68_0_2328_i_a7_0_0_a3_0_a3_0_a2_1_1_net_1), .C(
        Shift_reg_68_1_2300_i_0_o2), .D(\State1_ns_0_o5_2[0]_net_1 ), 
        .Y(Shift_reg_68_21_1723_i_i_a2_6_1_net_1));
    SLE \Parity_Counter[2]  (.D(\Parity_Counter_9[2]_net_1 ), .CLK(
        RX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Parity_Counter[2]_net_1 ));
    CFG3 #( .INIT(8'h04) )  Shift_reg_68_54_0 (.A(N_243), .B(
        Shift_reg_68_sn_N_49), .C(Shift_reg_68_sn_m37_u_i_0), .Y(
        Shift_reg_68_54_2));
    SLE \Shift_reg[1]  (.D(N_3652_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[1]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_14_1925_i_m4_ns (.A(
        Shift_reg_68_14_1925_i_m4_am_net_1), .B(
        Shift_reg_68_14_1925_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4417));
    CFG2 #( .INIT(4'h7) )  Shift_reg_68_28_12_1_i_o2_1 (.A(
        \State1[0]_net_1 ), .B(un14lto0), .Y(
        Shift_reg_68_28_12_1_i_o2_1_net_1));
    SLE \TC_Error_Counter[14]  (.D(\TC_Error_Counter_s[14] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[14]));
    CFG4 #( .INIT(16'h8008) )  Shift_reg_68_38_1263_i_a7_1_RNO (.A(
        \un1_Syn_reg[2] ), .B(N_53_i), .C(\un1_Syn_reg[0] ), .D(
        \un1_Syn_reg[6] ), .Y(N_1466));
    CFG4 #( .INIT(16'h0080) )  Shift_reg_68_28_28 (.A(
        \Bit_Counter[1]_net_1 ), .B(\Bit_Counter[2]_net_1 ), .C(
        Shift_reg_68_28_28_1_net_1), .D(N_86), .Y(
        Shift_reg_68_28_28_net_1));
    SLE \TC_Packet_Counter[5]  (.D(\TC_Packet_Counter_s[5] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[5]));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[37]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4226), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4223_i_0));
    CFG4 #( .INIT(16'h4544) )  Shift_reg_68_19_1783_i_0_1 (.A(
        Shift_reg_68_sn_N_84_mux), .B(
        Shift_reg_68_19_1783_i_0_a2_2_1_net_1), .C(
        \Shift_reg[34]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_19_1783_i_0_1_net_1));
    CFG3 #( .INIT(8'h40) )  Shift_reg_68_28_5_1 (.A(
        \Bit_Counter[1]_net_1 ), .B(\Bit_Counter[2]_net_1 ), .C(
        Shift_reg_68_28_6_4), .Y(Shift_reg_68_28_5_1_net_1));
    SLE \TC_Packet_Counter[24]  (.D(\TC_Packet_Counter_s[24] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[24]));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[2]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3630), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3627_i_0));
    CFG4 #( .INIT(16'hC080) )  \un1_Syn_reg_i_o3_RNIHOEC5[2]  (.A(
        Shift_reg_68_sn_m37_u_i_0), .B(\Shift_reg_68_54_e_0[11] ), .C(
        Shift_reg_68_sn_N_49), .D(N_243), .Y(N_1435));
    SLE \Parity_Counter[1]  (.D(\Parity_Counter_9[1]_net_1 ), .CLK(
        RX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Parity_Counter[1]_net_1 ));
    CFG4 #( .INIT(16'h0F53) )  DataO_10_iv_0_0_RNO_3 (.A(N_318), .B(
        N_2663), .C(\un22_DataO_i[1] ), .D(\un22_DataO_i[0] ), .Y(
        DataO_6_46_1_2));
    CFG4 #( .INIT(16'h0A0E) )  Flag_once_RNO (.A(
        un1_TC_Packet_Counter17_1_net_1), .B(N_2121), .C(N_2969_1), .D(
        un1_DataI), .Y(N_2969_i_0));
    CFG4 #( .INIT(16'h8000) )  TC_Packet_Counter18_i_a3 (.A(un14lto0), 
        .B(\Bit_Counter[1]_net_1 ), .C(N_21_i), .D(N_290), .Y(N_277));
    SLE \Shift_reg[55]  (.D(N_4464_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[55]_net_1 ));
    CFG2 #( .INIT(4'h4) )  Shift_reg_68_19_1783_i_0_a2_2_1 (.A(
        \un1_Syn_reg[6] ), .B(\un1_Syn_reg[0] ), .Y(N_417_1));
    SLE \Shift_reg[24]  (.D(N_3816_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[24]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  Shift_reg_68_6_2159_i_i_a2_3_2 (.A(
        \State1[0]_net_1 ), .B(TC_Packet_Counter17_i_0), .C(RX_GPIO0_c)
        , .D(CCA_NIRQ_c), .Y(Shift_reg_68_6_2159_i_i_a2_3_2_net_1));
    CFG4 #( .INIT(16'h0190) )  un1_Syn_reg_67_1_a2_0_0 (.A(
        \un1_Syn_reg[2] ), .B(\un1_Syn_reg[3]_net_1 ), .C(
        \un1_Syn_reg[6] ), .D(\un1_Syn_reg[5] ), .Y(r_m1_e_1));
    CFG4 #( .INIT(16'h9A00) )  Shift_reg_68_60_782_i_i_a2_0 (.A(
        \Shift_reg[9]_net_1 ), .B(Shift_reg_68_60_782_i_i_o2_2_0_net_1)
        , .C(Shift_reg_68_54_net_1), .D(N_250), .Y(N_193));
    CFG4 #( .INIT(16'h7F5F) )  un1_TC_Packet_Counter17_3 (.A(
        TC_Packet_Counter17_i_0), .B(
        un1_DataI_0_a3_a_a_a_a_a_a_N_5L7_net_1), .C(N_277), .D(
        un1_DataI_0_a3_a_a_a_a_a_a_x_net_1), .Y(
        un1_TC_Packet_Counter17_3_net_1));
    SLE \Parity[0]  (.D(N_3227_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_10_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Parity[0]_net_1 ));
    CFG4 #( .INIT(16'h3CF2) )  \un1_Syn_reg_RNIRK8I[3]  (.A(
        \un1_Syn_reg[3]_net_1 ), .B(\un1_Syn_reg[2] ), .C(N_53_i), .D(
        \un1_Syn_reg[6] ), .Y(Shift_reg_68_sn_N_42));
    CFG3 #( .INIT(8'h6A) )  Shift_reg_68_15_1897_i_m4_am (.A(
        \Shift_reg[30]_net_1 ), .B(\un1_Syn_reg[0] ), .C(N_1445), .Y(
        Shift_reg_68_15_1897_i_m4_am_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[9]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[9]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[8]_net_1 ), .S(
        \TC_Error_Counter_s[9] ), .Y(), .FCO(
        \TC_Error_Counter_cry[9]_net_1 ));
    CFG4 #( .INIT(16'h0C06) )  \Start_Sequence_counter_9[3]  (.A(
        SUM_m2_1), .B(\un6_DataO_i[3] ), .C(\un1_block_counter_7[0] ), 
        .D(SUM_m2_e), .Y(\Start_Sequence_counter_9[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  Shift_reg_68_28_0_0 (.A(
        \Bit_Counter[3]_net_1 ), .B(un14lto0), .C(N_385), .Y(
        Shift_reg_68_28_0_0_net_1));
    SLE \TC_Packet_Counter[23]  (.D(\TC_Packet_Counter_s[23] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[23]));
    CFG2 #( .INIT(4'h1) )  \Parity_Counter_9[0]  (.A(
        \un1_block_counter_4[0]_net_1 ), .B(N_143), .Y(
        \Parity_Counter_9[0]_net_1 ));
    CFG4 #( .INIT(16'h4C44) )  Block_ErrO_2_sqmuxa_1_i_a0_0_RNIP1OP3 (
        .A(TC_Packet_Counter17_i_0), .B(Block_ErrO_2_sqmuxa_1_i_a1_0), 
        .C(un1_TC_Packet_Counter17_3_net_1), .D(Shift_N_7_1), .Y(
        N_79_i_1));
    SLE \Bit_Counter[3]  (.D(\Bit_Counter_lm[3] ), .CLK(RX_GPIO1_c), 
        .EN(un1_DataO41_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Bit_Counter[3]_net_1 ));
    SLE \Parity[6]  (.D(N_3700_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_10_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Parity[6]_net_1 ));
    CFG4 #( .INIT(16'hFEBA) )  \un1_Syn_reg_i_o3_0_x2_RNIDEP63[1]  (.A(
        N_53_i), .B(N_1431), .C(Shift_reg_68_sn_m72_6_am_1), .D(
        Shift_reg_68_sn_m59_i_x3_RNI590H_net_1), .Y(
        \un1_Syn_reg_i_o3_0_x2_RNIDEP63[1]_net_1 ));
    SLE \Start_Buff[13]  (.D(N_3366), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[13]_net_1 ));
    CFG3 #( .INIT(8'hFD) )  Shift_reg_68_9_2070_i_0_o2_1_1 (.A(
        \Bit_Counter[1]_net_1 ), .B(un14lto4), .C(N_55), .Y(
        Shift_reg_68_9_2070_i_0_o2_1_1_net_1));
    CFG4 #( .INIT(16'h4F7F) )  Shift_reg_68_57_866_i_i_0_RNO_0 (.A(
        N_90), .B(N_82), .C(\Shift_reg[6]_net_1 ), .D(N_123), .Y(
        Shift_reg_68_57_866_i_i_0_RNO_0_net_1));
    CFG3 #( .INIT(8'h82) )  DataO_0_sqmuxa_1_0 (.A(CCA_NIRQ_c), .B(
        \State2[0]_net_1 ), .C(\State2[1]_net_1 ), .Y(
        DataO_0_sqmuxa_1_0_net_1));
    CFG2 #( .INIT(4'h7) )  Shift_reg_68_28_1_0_o2 (.A(
        \Bit_Counter[3]_net_1 ), .B(\Bit_Counter[1]_net_1 ), .Y(N_91));
    CFG4 #( .INIT(16'h1131) )  Shift_reg_68_39_1233_i_a7 (.A(
        \State1[0]_net_1 ), .B(\Shift_reg[23]_net_1 ), .C(
        Shift_reg_68_sn_N_73), .D(un1_TC_Packet_Counter17_3_net_1), .Y(
        N_3842));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[7]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3511), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3508_i_0));
    SLE \Start_Sequence_counter[2]  (.D(
        \Start_Sequence_counter_9[2]_net_1 ), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\un6_DataO_i[2] ));
    CFG2 #( .INIT(4'h8) )  \Bit_Counter_lm_0[5]  (.A(
        Bit_Counter_3_sqmuxa), .B(\Bit_Counter_s[5]_net_1 ), .Y(
        \Bit_Counter_lm[5] ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[11]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[11]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[10]_net_1 ), .S(
        \TC_Error_Counter_s[11] ), .Y(), .FCO(
        \TC_Error_Counter_cry[11]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \Shift_reg_RNIU5E6[27]  (.A(
        \Shift_reg[27]_net_1 ), .B(\Shift_reg[25]_net_1 ), .C(
        \Shift_reg[19]_net_1 ), .D(\Shift_reg[13]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_43));
    CFG2 #( .INIT(4'h8) )  Shift_reg_68_28_12_0 (.A(N_436_1), .B(
        Shift_reg_68_28_9_2), .Y(Shift_reg_68_28_12_0_net_1));
    CFG2 #( .INIT(4'h7) )  Parity_16_1_505_i_0_o2_0 (.A(
        \Parity_Counter[1]_net_1 ), .B(\Parity_Counter[2]_net_1 ), .Y(
        Parity_16_1_505_i_0_o2_0_net_1));
    CFG4 #( .INIT(16'h1468) )  Shift_reg_68_sn_m57_1_RNIVNOR_0 (.A(
        \un1_Syn_reg[2] ), .B(\un1_Syn_reg[5] ), .C(\un1_Syn_reg[4] ), 
        .D(\un1_Syn_reg[3]_net_1 ), .Y(Shift_reg_68_sn_m72_6_am_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[25]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[25]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[24]_net_1 ), .S(
        \TC_Error_Counter_s[25] ), .Y(), .FCO(
        \TC_Error_Counter_cry[25]_net_1 ));
    SLE \Shift_reg[8]  (.D(N_3483_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[8]_net_1 ));
    CFG4 #( .INIT(16'hFCF5) )  Shift_reg_68_20_1753_i_2 (.A(
        \Shift_reg[35]_net_1 ), .B(Shift_reg_68_20_1753_i_a7_1_0_net_1)
        , .C(Shift_reg_68_20_1753_i_0_net_1), .D(
        Shift_reg_68_sn_N_84_mux), .Y(Shift_reg_68_20_1753_i_2_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[29]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[29]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[28]_net_1 ), .S(
        \TC_Error_Counter_s[29] ), .Y(), .FCO(
        \TC_Error_Counter_cry[29]_net_1 ));
    SLE \TC_Error_Counter[4]  (.D(\TC_Error_Counter_s[4] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[4]));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_59_810_i_m4_ns (.A(
        Shift_reg_68_59_810_i_m4_am_net_1), .B(
        Shift_reg_68_59_810_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3486));
    ARI1 #( .INIT(20'h40800) )  \Shift_Bit_Counter_cry_cy[0]  (.A(
        N_302), .B(CCA_NIRQ_c), .C(\State2[0]_net_1 ), .D(
        \State2[1]_net_1 ), .FCI(VCC_net_1), .S(), .Y(
        \Shift_Bit_Counter_cry_cy_Y[0] ), .FCO(
        Shift_Bit_Counter_cry_cy));
    SLE DataO (.D(DataO_10), .CLK(RX_GPIO1_c), .EN(un1_DataO41_14_i_0), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(A_1));
    CFG4 #( .INIT(16'hFFDF) )  Shift_reg_68_23_1667_i_i_o3 (.A(
        Shift_reg_68_28_30_3), .B(N_87), .C(un14lto4), .D(un14lto5), 
        .Y(N_216));
    CFG4 #( .INIT(16'h0008) )  un1_DataI_0_a3_a_a_a_a_a_a_N_2L1 (.A(
        \Shift_reg[46]_net_1 ), .B(\Shift_reg[40]_net_1 ), .C(
        \Shift_reg[9]_net_1 ), .D(\Shift_reg[4]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_N_2L1_net_1));
    CFG3 #( .INIT(8'h04) )  Shift_reg_68_28_1_1 (.A(
        \Bit_Counter[1]_net_1 ), .B(\Bit_Counter[3]_net_1 ), .C(N_385), 
        .Y(Shift_reg_68_28_1_1_net_1));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_28_3_a2_0_a3 (.A(
        \Bit_Counter[3]_net_1 ), .B(un14lto4), .C(un14lto5), .Y(
        Shift_reg_68_28_6_4));
    CFG4 #( .INIT(16'hFFFE) )  \State1_ns_0_o5_3[0]  (.A(un1_Syn_reg_2)
        , .B(N_2847), .C(N_2846), .D(N_2843), .Y(
        \State1_ns_0_o5_3[0]_net_1 ));
    CFG4 #( .INIT(16'h0405) )  \Shift_reg_RNO[34]  (.A(
        Shift_reg_68_19_1783_i_0_0_net_1), .B(\Shift_reg[34]_net_1 ), 
        .C(Shift_reg_68_19_1783_i_0_1_net_1), .D(N_388), .Y(N_4292_i_0)
        );
    CFG4 #( .INIT(16'h0004) )  un1_Syn_reg_2_0_a3_RNI6MOJ1 (.A(
        un1_Syn_reg_2), .B(\State1[0]_net_1 ), .C(N_2846), .D(N_2847), 
        .Y(un1_Syn_reg_2_0_a3_RNI6MOJ1_net_1));
    CFG4 #( .INIT(16'h0001) )  un1_Start_Buff_1_11 (.A(
        \Start_Buff[3]_net_1 ), .B(\Start_Buff[2]_net_1 ), .C(
        \Start_Buff[1]_net_1 ), .D(\Start_Buff[0]_net_1 ), .Y(
        un1_Start_Buff_1_11_net_1));
    CFG2 #( .INIT(4'h1) )  Shift_reg_68_43_1_0_a2 (.A(\un1_Syn_reg[0] )
        , .B(\un1_Syn_reg[5] ), .Y(Shift_reg_68_43_2));
    CFG4 #( .INIT(16'h78F0) )  Shift_reg_68_32_1435_i_m4_am (.A(
        \Shift_reg_68_54_e_0[8] ), .B(Shift_reg_68_54_2), .C(
        \Shift_reg[16]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_32_1435_i_m4_am_net_1));
    CFG4 #( .INIT(16'hF0B8) )  Parity_16_1089_i_m5 (.A(RX_GPIO0_c), .B(
        \Parity_Counter[0]_net_1 ), .C(\Parity[5]_net_1 ), .D(N_3721), 
        .Y(N_3723));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIL6T18[26]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[26]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[25] ), .S(
        \TC_Packet_Counter_s[26] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[26] ));
    SLE \Shift_reg[39]  (.D(N_4176_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[39]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_18_1811_i_m4_ns (.A(
        Shift_reg_68_18_1811_i_m4_am_net_1), .B(
        Shift_reg_68_18_1811_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4320));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[48]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4630), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4627_i_0));
    CFG3 #( .INIT(8'hFD) )  Shift_reg_68_1_2300_i_0_o3_0 (.A(
        Shift_reg_68_sn_N_49), .B(Shift_reg_68_1_2300_i_0_o3_0_0_net_1)
        , .C(Shift_reg_68_sn_m37_u_i_0), .Y(N_392));
    CFG2 #( .INIT(4'h8) )  Shift_reg_68_28_21_i_a2_1 (.A(
        \Bit_Counter[2]_net_1 ), .B(\Bit_Counter[3]_net_1 ), .Y(N_290));
    CFG2 #( .INIT(4'h1) )  Shift_reg_68_13_1953_i_i_N_4L5_N_4L6 (.A(
        N_90), .B(N_91), .Y(Shift_reg_68_13_1953_i_i_N_4L5_N_4L6_net_1)
        );
    CFG2 #( .INIT(4'h8) )  Shift_reg_68_42_1143_i_m4_am_RNO (.A(
        Shift_reg_68_sn_N_16), .B(\un1_Syn_reg[5] ), .Y(
        \Shift_reg_68_54_e_0[26] ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[16]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[16]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[15]_net_1 ), .S(
        \TC_Error_Counter_s[16] ), .Y(), .FCO(
        \TC_Error_Counter_cry[16]_net_1 ));
    SLE \Syn_reg[2]  (.D(N_3301_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_15_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Syn_reg[2]_net_1 ));
    CFG4 #( .INIT(16'hA0DD) )  DataO_10_iv_0_a3_0_RNO (.A(
        \un6_DataO_i[0] ), .B(N_2627), .C(N_2624), .D(DataO_2_15_1_2), 
        .Y(DataO_2));
    CFG4 #( .INIT(16'hE800) )  un1_DataO41_22_0_a2_0 (.A(
        \un1_Syn_reg[5] ), .B(\un1_Syn_reg[6] ), .C(
        \un1_Syn_reg[3]_net_1 ), .D(N_370), .Y(N_373));
    SLE \Shift_reg[14]  (.D(N_67), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[14]_net_1 ));
    CFG3 #( .INIT(8'h14) )  \Syn_reg_RNO[0]  (.A(N_54), .B(RX_GPIO0_c), 
        .C(\Syn_reg[6]_net_1 ), .Y(N_3332_i_0));
    SLE \Shift_reg[25]  (.D(N_3792_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[25]_net_1 ));
    CFG4 #( .INIT(16'hFD20) )  Parity_16_2_480_i_0_m2 (.A(
        \Parity_Counter[0]_net_1 ), .B(Parity_16_3_456_i_o4_0), .C(
        RX_GPIO0_c), .D(\Parity[1]_net_1 ), .Y(N_80));
    CFG4 #( .INIT(16'h0109) )  \Shift_reg_RNO_0[44]  (.A(
        \un1_Syn_reg[0] ), .B(\Shift_reg[44]_net_1 ), .C(
        Shift_reg_68_sn_N_84_mux), .D(N_392), .Y(N_4727_i_1));
    ARI1 #( .INIT(20'h48800) )  \Shift_Bit_Counter_cry[4]  (.A(
        VCC_net_1), .B(\Shift_Bit_Counter[4]_net_1 ), .C(
        \Shift_Bit_Counter_cry_cy_Y[0] ), .D(GND_net_1), .FCI(
        \Shift_Bit_Counter_cry[3]_net_1 ), .S(\Shift_Bit_Counter_s[4] )
        , .Y(), .FCO(\Shift_Bit_Counter_cry[4]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_27_1552_i_m4_ns (.A(
        Shift_reg_68_27_1552_i_m4_am_net_1), .B(
        Shift_reg_68_27_1552_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4104));
    CFG2 #( .INIT(4'h8) )  \un1_Syn_reg_i_o3_RNIETLE4[2]  (.A(
        Shift_reg_68_sn_N_49), .B(\Shift_reg_68_54_e_0[42] ), .Y(
        N_1461));
    CFG4 #( .INIT(16'h0800) )  Shift_reg_68_60_782_i_i_0_RNO (.A(
        \Shift_reg[9]_net_1 ), .B(\State1[0]_net_1 ), .C(
        Shift_reg_68_1_2300_i_0_o2), .D(N_220), .Y(Shift_m3_0_a2_2_2));
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_2_2272_i_m4_bm (.A(
        Shift_reg_68_28_0_0_net_1), .B(N_374), .C(RX_GPIO0_c), .D(
        \Shift_reg[45]_net_1 ), .Y(Shift_reg_68_2_2272_i_m4_bm_net_1));
    CFG4 #( .INIT(16'h0040) )  un1_Syn_reg_67_1_a2_0_0_RNIN2II1 (.A(
        \un1_Syn_reg[0] ), .B(r_m1_e_1), .C(\un1_Syn_reg[4] ), .D(
        N_53_i), .Y(N_2843));
    CFG4 #( .INIT(16'h0F8F) )  Shift_reg_68_63_697_i_i_1 (.A(
        Shift_reg_68_63_697_i_i_a2_3_0_net_1), .B(Shift_m2_1_1), .C(
        Shift_reg_68_63_697_i_i_N_5L8_net_1), .D(Shift_N_5), .Y(
        Shift_reg_68_63_697_i_i_1_0));
    CFG4 #( .INIT(16'h0C06) )  \Start_Sequence_counter_9[1]  (.A(
        \un6_DataO_i[0] ), .B(\un6_DataO_i[1] ), .C(
        \un1_block_counter_7[0] ), .D(un1_DataO41_18), .Y(
        \Start_Sequence_counter_9[1]_net_1 ));
    SLE \Shift_reg[32]  (.D(N_4342_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[32]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIUIRD2[3]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[3]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Packet_Counter_cry[2] ), .S(
        \TC_Packet_Counter_s[3] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[3] ));
    SLE \Start_Sequence_counter[0]  (.D(
        \Start_Sequence_counter_9[0]_net_1 ), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\un6_DataO_i[0] ));
    SLE \Shift_reg[53]  (.D(N_4511_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[53]_net_1 ));
    CFG3 #( .INIT(8'h04) )  Shift_reg_68_57_866_i_i_RNO (.A(N_90), .B(
        N_253), .C(N_102), .Y(Shift_N_10_mux));
    CFG4 #( .INIT(16'h0080) )  \Parity_RNO[6]  (.A(CCA_NIRQ_c), .B(
        TC_Packet_Counter17_i_0), .C(N_3703), .D(N_277), .Y(N_3700_i_0)
        );
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNII5N26[15]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[15]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[14] ), .S(
        \TC_Packet_Counter_s[15] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[15] ));
    SLE \Start_Buff[2]  (.D(N_3112), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[2]_net_1 ));
    CFG4 #( .INIT(16'h530F) )  DataO_10_iv_0_a3_0_RNO_8 (.A(
        \Start_Buff[3]_net_1 ), .B(\Start_Buff[7]_net_1 ), .C(
        \un6_DataO_i[2] ), .D(\un6_DataO_i[3] ), .Y(DataO_2_3_1_2));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_9_2070_i_0_a3_0 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(
        Shift_reg_68_9_2070_i_0_a3_0_0_net_1), .D(N_82), .Y(N_285));
    CFG3 #( .INIT(8'h04) )  Shift_reg_68_21_1723_i_i_3_RNO (.A(N_90), 
        .B(N_253), .C(N_100), .Y(N_227));
    SLE \Start_Buff[0]  (.D(N_3132), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[0]_net_1 ));
    CFG4 #( .INIT(16'h3020) )  Shift_reg_68_sn_m57_i_o3_RNIR79Q (.A(
        \un1_Syn_reg[5] ), .B(N_53_i), .C(\un1_Syn_reg[0] ), .D(
        \un1_Syn_reg[6] ), .Y(N_243));
    CFG4 #( .INIT(16'h195D) )  DataO_10_iv_0_0_RNO_10 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[8]_net_1 ), .D(\Shift_reg[12]_net_1 ), .Y(
        DataO_6_44_1_2));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[54]  (.A(
        Shift_reg_68_28_9_0_net_1), .B(N_86), .C(RX_GPIO0_c), .D(
        \Shift_reg[54]_net_1 ), .Y(N_124));
    CFG4 #( .INIT(16'hF3F7) )  Shift_reg_68_19_1783_i_0_o3_0 (.A(N_243)
        , .B(Shift_reg_68_sn_N_49), .C(N_97_i), .D(
        Shift_reg_68_sn_m37_u_i_0), .Y(N_381));
    CFG4 #( .INIT(16'h0010) )  Shift_reg_68_30_1493_i_i_0_RNO_1 (.A(
        \un1_Syn_reg[5] ), .B(\Shift_reg[14]_net_1 ), .C(
        \un1_Syn_reg[6] ), .D(N_53_i), .Y(Shift_m2_0_0));
    ARI1 #( .INIT(20'h48800) )  \Shift_Bit_Counter_cry[2]  (.A(
        VCC_net_1), .B(\un22_DataO_i[2] ), .C(
        \Shift_Bit_Counter_cry_cy_Y[0] ), .D(GND_net_1), .FCI(
        \Shift_Bit_Counter_cry[1]_net_1 ), .S(\Shift_Bit_Counter_s[2] )
        , .Y(), .FCO(\Shift_Bit_Counter_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIIHKG7[23]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[23]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[22] ), .S(
        \TC_Packet_Counter_s[23] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[23] ));
    CFG4 #( .INIT(16'hAAA2) )  un1_TC_Packet_Counter17_3_RNIHKFMA (.A(
        \State1[0]_net_1 ), .B(
        \un1_Syn_reg_i_o3_0_x2_RNIDEP63[1]_net_1 ), .C(
        Shift_reg_68_sn_m72_7_ns_sx), .D(
        un1_TC_Packet_Counter17_3_net_1), .Y(Shift_reg_68_sn_N_84_mux));
    CFG4 #( .INIT(16'h0040) )  \un1_Syn_reg_i_o3_0_x2_RNIV1AC5[1]  (.A(
        Shift_reg_68_sn_m37_u_i_0), .B(\Shift_reg_68_54_e_0[30] ), .C(
        Shift_reg_68_sn_N_49), .D(N_243), .Y(N_1445));
    CFG4 #( .INIT(16'hEAAA) )  un1_DataO41_22_0_0 (.A(un1_CCA_i_0), .B(
        Bit_Counter_3_sqmuxa), .C(\Bit_Counter[3]_net_1 ), .D(N_21_i), 
        .Y(un1_DataO41_22_0_0_net_1));
    CFG4 #( .INIT(16'h3F15) )  \Shift_reg_RNO_0[32]  (.A(N_349_1), .B(
        un1_TC_Packet_Counter17_5_net_1), .C(\State1[0]_net_1 ), .D(
        N_1452_mux), .Y(N_4342_i_1));
    CFG4 #( .INIT(16'hEDCC) )  Shift_reg_68_46_1115_i_i (.A(
        Shift_reg_68_46_1115_i_i_N_7L14_net_1), .B(
        Shift_reg_68_46_1115_i_i_1), .C(\Shift_reg[27]_net_1 ), .D(
        N_250), .Y(N_69));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[10]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[10]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[9]_net_1 ), .S(
        \TC_Error_Counter_s[10] ), .Y(), .FCO(
        \TC_Error_Counter_cry[10]_net_1 ));
    CFG2 #( .INIT(4'h4) )  Shift_reg_68_9_2070_i_0_a3_0_0 (.A(N_268), 
        .B(\Shift_reg[52]_net_1 ), .Y(
        Shift_reg_68_9_2070_i_0_a3_0_0_net_1));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[51]  (.A(
        Shift_reg_68_28_6_0_net_1), .B(N_92), .C(RX_GPIO0_c), .D(
        \Shift_reg[51]_net_1 ), .Y(N_121));
    CFG4 #( .INIT(16'h0C26) )  Shift_reg_68_26_1580_i_i_N_7L13 (.A(
        Shift_reg_68_26_1580_i_i_1_tz_net_1), .B(\Shift_reg[41]_net_1 )
        , .C(Shift_reg_68_13_1953_i_i_o3_0_0_net_1), .D(N_74), .Y(
        Shift_reg_68_26_1580_i_i_1));
    CFG4 #( .INIT(16'hF780) )  Shift_reg_68_47_1039_i_m4_0_bm (.A(
        N_21_i), .B(Shift_reg_68_28_3_4), .C(RX_GPIO0_c), .D(
        \Shift_reg[0]_net_1 ), .Y(Shift_reg_68_47_1039_i_m4_0_bm_net_1)
        );
    CFG4 #( .INIT(16'h0D05) )  Shift_reg_1_sqmuxa_1_i_o3_0_o2_RNIHTIS 
        (.A(CCA_NIRQ_c), .B(\State1[0]_net_1 ), .C(un1_CCA_i_0), .D(
        N_58), .Y(un1_DataO41_10_i_0));
    CFG2 #( .INIT(4'h6) )  Shift_reg_68_sn_m57_1 (.A(\Parity[4]_net_1 )
        , .B(\Syn_reg[4]_net_1 ), .Y(\un1_Syn_reg[4] ));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_0_668_a2 (.A(CCA_NIRQ_c), .B(
        \Start_Buff[13]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3356));
    CFG4 #( .INIT(16'hFFFB) )  Shift_reg_68_46_1115_i_i_o3 (.A(
        un14lto0), .B(\Bit_Counter[3]_net_1 ), .C(N_92), .D(N_110), .Y(
        N_215));
    CFG4 #( .INIT(16'h9621) )  \State1_ns_0_o5_2[0]  (.A(
        \un1_Syn_reg[0] ), .B(N_73_i), .C(\un1_Syn_reg[4] ), .D(N_53_i)
        , .Y(\State1_ns_0_o5_2[0]_net_1 ));
    CFG4 #( .INIT(16'hFFF4) )  Shift_reg_68_63_697_i_i (.A(
        Shift_reg_68_1_2300_i_0_o2_0_RNIHMNKG_net_1), .B(
        \Shift_reg[12]_net_1 ), .C(N_199_1), .D(
        Shift_reg_68_63_697_i_i_1_0), .Y(N_75));
    CFG4 #( .INIT(16'hF5F7) )  Shift_reg_68_31_1463_i_1 (.A(CCA_NIRQ_c)
        , .B(\Shift_reg[15]_net_1 ), .C(N_4036), .D(
        Shift_reg_68_sn_N_84_mux), .Y(Shift_reg_68_31_1463_i_1_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \Bit_Counter_cry[3]  (.A(VCC_net_1), 
        .B(\Bit_Counter[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \Bit_Counter_cry[2]_net_1 ), .S(\Bit_Counter_s[3] ), .Y(), 
        .FCO(\Bit_Counter_cry[3]_net_1 ));
    CFG4 #( .INIT(16'hFF37) )  Shift_reg_68_8_2099_i_0_1 (.A(
        \Shift_reg[51]_net_1 ), .B(CCA_NIRQ_c), .C(
        Shift_reg_68_sn_N_84_mux), .D(N_350), .Y(
        Shift_reg_68_8_2099_i_0_1_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[8]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[8]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[7]_net_1 ), .S(
        \TC_Error_Counter_s[8] ), .Y(), .FCO(
        \TC_Error_Counter_cry[8]_net_1 ));
    SLE \TC_Error_Counter[23]  (.D(\TC_Error_Counter_s[23] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[23]));
    CFG3 #( .INIT(8'h04) )  \Shift_reg_RNO[5]  (.A(
        Shift_reg_68_56_895_i_1_net_1), .B(N_3558_i_1), .C(N_3563), .Y(
        N_3558_i_0));
    CFG3 #( .INIT(8'h04) )  \Shift_reg_RNO[32]  (.A(
        Shift_reg_68_17_1839_i_1_net_1), .B(N_4342_i_1), .C(N_4347), 
        .Y(N_4342_i_0));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h2) )  un1_DataO41_24_i_a3_1 (.A(
        un1_block_counter_net_1), .B(CCA_NIRQ_c), .Y(N_357));
    CFG3 #( .INIT(8'h04) )  \Shift_reg_RNO[15]  (.A(
        Shift_reg_68_31_1463_i_1_net_1), .B(N_4032_i_1), .C(N_4037), 
        .Y(N_4032_i_0));
    SLE \Shift_reg[44]  (.D(N_4727_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[44]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIJS8N5[13]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[13]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[12] ), .S(
        \TC_Packet_Counter_s[13] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[13] ));
    CFG4 #( .INIT(16'hAAEA) )  Shift_reg_68_19_1783_i_0_0 (.A(N_74), 
        .B(Shift_reg_68_sn_N_84_mux), .C(N_287), .D(N_104), .Y(
        Shift_reg_68_19_1783_i_0_0_net_1));
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_62_726_i_m4_bm (.A(
        Shift_reg_68_28_51_0_net_1), .B(N_92), .C(RX_GPIO0_c), .D(
        \Shift_reg[11]_net_1 ), .Y(Shift_reg_68_62_726_i_m4_bm_net_1));
    CFG4 #( .INIT(16'h0020) )  Shift_reg_68_30_1493_i_i_0_RNO_0 (.A(
        Shift_reg_1_sqmuxa_1_i_o3_0_o2_RNIJK1N_0_net_1), .B(
        Shift_reg_68_sn_N_56), .C(Shift_m2_0_0), .D(
        Shift_reg_68_1_2300_i_0_o2), .Y(Shift_m2_0_3));
    CFG4 #( .INIT(16'hFFF4) )  Shift_reg_68_60_782_i_i (.A(N_220), .B(
        N_253), .C(Shift_reg_68_60_782_i_i_0_net_1), .D(N_193), .Y(
        N_73));
    CFG4 #( .INIT(16'h13FF) )  un1_DataO41_18_1 (.A(N_152), .B(
        TC_Packet_Counter18_i_0), .C(N_356_1), .D(N_3002), .Y(
        un1_DataO41_18_1_net_1));
    SLE \Shift_reg[15]  (.D(N_4032_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[15]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  Shift_reg_68_28_18_a2_0_o2 (.A(
        \Bit_Counter[2]_net_1 ), .B(un14lto5), .C(
        \Bit_Counter[3]_net_1 ), .Y(N_55));
    CFG4 #( .INIT(16'h8000) )  un1_Syn_reg_2_0_a3 (.A(N_244_2), .B(
        \un1_Syn_reg[3]_net_1 ), .C(N_370), .D(N_94_i), .Y(
        un1_Syn_reg_2));
    CFG4 #( .INIT(16'h5955) )  \Parity_Counter_9_RNO[0]  (.A(
        \Parity_Counter[0]_net_1 ), .B(\State1[0]_net_1 ), .C(
        un1_CCA_i_0), .D(N_58), .Y(N_143));
    SLE \Shift_reg[36]  (.D(N_56), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[36]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  Shift_reg_68_1_2300_i_0_o2_0_RNIHMNKG (.A(
        un1_TC_Packet_Counter17_3_RNIS3QPC_net_1), .B(
        Shift_reg_68_1_2300_i_0_o2), .C(Shift_N_7_mux_2), .Y(
        Shift_reg_68_1_2300_i_0_o2_0_RNIHMNKG_net_1));
    CFG3 #( .INIT(8'hAC) )  \un1_Syn_reg_i_o3_RNITFTS6[6]  (.A(
        Shift_reg_68_sn_m59_i_x3_RNI3Q7P3_net_1), .B(
        Shift_reg_68_sn_m72_6_ns_1), .C(\un1_Syn_reg[6] ), .Y(N_2551));
    SLE \Shift_reg[23]  (.D(N_3841_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[23]_net_1 ));
    CFG3 #( .INIT(8'h12) )  \block_counter_8[1]  (.A(CO0), .B(
        \un1_block_counter_7[0] ), .C(\block_counter[1]_net_1 ), .Y(
        \block_counter_8[1]_net_1 ));
    SLE \TC_Error_Counter[10]  (.D(\TC_Error_Counter_s[10] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[10]));
    CFG4 #( .INIT(16'h00B3) )  Shift_reg_68_12_1982_i_m4_am_RNO_0 (.A(
        \un1_Syn_reg[0] ), .B(\State1[0]_net_1 ), .C(
        Shift_reg_68_sn_N_32), .D(Shift_reg_68_sn_N_78_mux), .Y(
        \Shift_reg_68_54_e_1[55] ));
    CFG4 #( .INIT(16'h6006) )  \Syn_reg_RNI2RFH1[1]  (.A(
        \Parity[1]_net_1 ), .B(\Syn_reg[1]_net_1 ), .C(
        \Syn_reg[6]_net_1 ), .D(\Parity[6]_net_1 ), .Y(
        \Syn_reg_RNI2RFH1[1]_net_1 ));
    SLE \Shift_reg[38]  (.D(N_63), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[38]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \Shift_reg_RNIFPPJ1[10]  (.A(
        un1_DataI_0_a3_a_a_a_a_a_a_0_36), .B(
        un1_DataI_0_a3_a_a_a_a_a_a_0_38), .C(
        un1_DataI_0_a3_a_a_a_a_a_a_0_37), .D(
        un1_DataI_0_a3_a_a_a_a_a_a_0_35), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_56));
    CFG4 #( .INIT(16'h0080) )  \Parity_RNO[4]  (.A(CCA_NIRQ_c), .B(
        TC_Packet_Counter17_i_0), .C(N_3150), .D(N_277), .Y(N_3147_i_0)
        );
    CFG4 #( .INIT(16'hECCC) )  DataO15_0_o2 (.A(\Bit_Counter[1]_net_1 )
        , .B(un14lto4), .C(un14lto0), .D(N_290), .Y(N_152));
    CFG3 #( .INIT(8'hBF) )  Shift_reg_68_6_2159_i_i_o2_0 (.A(
        \un1_Syn_reg[0] ), .B(Shift_reg_68_sn_m37_u_i_0), .C(
        Shift_reg_68_sn_N_49), .Y(N_101));
    CFG4 #( .INIT(16'h9030) )  Shift_reg_68_38_1263_i_a7_1 (.A(
        \un1_Syn_reg[0] ), .B(\Shift_reg[22]_net_1 ), .C(N_349_1), .D(
        N_1466), .Y(N_3866));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[10]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3436), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3433_i_0));
    CFG4 #( .INIT(16'hEB97) )  Shift_reg_68_sn_m57_1_RNIVNOR (.A(
        \un1_Syn_reg[2] ), .B(\un1_Syn_reg[5] ), .C(\un1_Syn_reg[4] ), 
        .D(\un1_Syn_reg[3]_net_1 ), .Y(N_41));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_0_2328_i_a7_2 (.A(
        Shift_reg_68_sn_N_56), .B(\Shift_reg[43]_net_1 ), .C(N_82), .Y(
        N_4756));
    CFG4 #( .INIT(16'h1230) )  \Parity_Counter_9[2]  (.A(CO0_0), .B(
        \un1_block_counter_4[0]_net_1 ), .C(\Parity_Counter[2]_net_1 ), 
        .D(\Parity_Counter[1]_net_1 ), .Y(\Parity_Counter_9[2]_net_1 ));
    CFG4 #( .INIT(16'h007F) )  un1_DataO41_27_a0_0_RNIMPF32 (.A(
        un1_DataO41_27_a0_0_net_1), .B(Syn_reg_0_sqmuxa_2_net_1), .C(
        N_2121), .D(un1_DataO41_1), .Y(un1_DataO41_27_i_0));
    CFG4 #( .INIT(16'hF078) )  Shift_reg_68_33_1407_i_m4_am (.A(
        \Shift_reg_68_54_e_0[17] ), .B(Shift_reg_68_54_net_1), .C(
        \Shift_reg[17]_net_1 ), .D(N_53_i), .Y(
        Shift_reg_68_33_1407_i_m4_am_net_1));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_29_1522_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_82), 
        .D(N_83), .Y(N_4084));
    SLE \TC_Packet_Counter[22]  (.D(\TC_Packet_Counter_s[22] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[22]));
    CFG4 #( .INIT(16'h9CCC) )  Shift_reg_68_22_1695_i_m4_am (.A(N_53_i)
        , .B(\Shift_reg[37]_net_1 ), .C(Shift_reg_68_54_2), .D(N_417_1)
        , .Y(Shift_reg_68_22_1695_i_m4_am_net_1));
    CFG3 #( .INIT(8'h15) )  Syn_reg_0_sqmuxa_0_RNI93JH (.A(un1_CCA_i_0)
        , .B(Syn_reg_0_sqmuxa_2_net_1), .C(Syn_reg_0_sqmuxa_0_net_1), 
        .Y(un1_DataO41_15_i_0));
    CFG4 #( .INIT(16'h78F0) )  Shift_reg_68_55_925_i_m4_am (.A(
        \Shift_reg_68_54_e_0[4] ), .B(Shift_reg_68_54_net_1), .C(
        \Shift_reg[4]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_55_925_i_m4_am_net_1));
    CFG4 #( .INIT(16'hF780) )  \Shift_reg_68_28[32]  (.A(
        Shift_reg_68_28_14_1), .B(Shift_reg_68_28_3_4), .C(RX_GPIO0_c), 
        .D(\Shift_reg[32]_net_1 ), .Y(N_102_0));
    CFG4 #( .INIT(16'hEFAA) )  Shift_reg_68_37_1293_i_0_1 (.A(N_74), 
        .B(Shift_reg_68_sn_N_84_mux), .C(N_402), .D(
        Shift_reg_68_37_1293_i_0_1_1_net_1), .Y(
        Shift_reg_68_37_1293_i_0_1_net_1));
    CFG2 #( .INIT(4'h4) )  Shift_reg_68_28_32_0 (.A(N_387), .B(
        Shift_reg_68_28_32_2_net_1), .Y(Shift_reg_68_28_32_0_net_1));
    CFG3 #( .INIT(8'h10) )  Shift_reg_68_54_11 (.A(
        Shift_reg_68_sn_N_32), .B(Shift_reg_68_sn_N_49), .C(
        \State1[0]_net_1 ), .Y(Shift_reg_68_54_4));
    CFG4 #( .INIT(16'h8000) )  un1_DataO41_24_i_a3_0_4 (.A(
        un1_DataO41_24_i_a3_0_1_net_1), .B(N_356_1), .C(N_3002), .D(
        N_152), .Y(un1_DataO41_24_i_a3_0_4_net_1));
    CFG3 #( .INIT(8'hAC) )  \un1_Syn_reg_RNIN54G2[3]  (.A(
        \un1_Syn_reg_RNIQLBC[3]_net_1 ), .B(Shift_reg_68_sn_m47_0_ns_1)
        , .C(\Syn_reg_RNI2RFH1[1]_net_1 ), .Y(N_2176));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_63_697_i_i_a2_3_0 (.A(
        \Shift_reg[12]_net_1 ), .B(Shift_reg_68_sn_N_9), .C(
        \un1_Syn_reg[5] ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_63_697_i_i_a2_3_0_net_1));
    CFG4 #( .INIT(16'h2000) )  \un1_Start_Sequence_counter_1.SUM_m2_1  
        (.A(\un6_DataO_i[2] ), .B(un1_DataO41_18_1_net_1), .C(
        \un6_DataO_i[1] ), .D(\un6_DataO_i[0] ), .Y(SUM_m2_1));
    SLE \TC_Error_Counter[6]  (.D(\TC_Error_Counter_s[6] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[6]));
    SLE \Start_Sequence_counter[3]  (.D(
        \Start_Sequence_counter_9[3]_net_1 ), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\un6_DataO_i[3] ));
    SLE \TC_Packet_Counter[7]  (.D(\TC_Packet_Counter_s[7] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[7]));
    SLE \TC_Packet_Counter[16]  (.D(\TC_Packet_Counter_s[16] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[16]));
    SLE \Start_Buff[5]  (.D(N_3082), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[5]_net_1 ));
    CFG4 #( .INIT(16'h1248) )  un1_Syn_reg_2_0_a3_1 (.A(
        \Syn_reg[1]_net_1 ), .B(\Syn_reg[0]_net_1 ), .C(
        \Parity[1]_net_1 ), .D(\Parity[0]_net_1 ), .Y(N_244_2));
    SLE \Shift_reg[45]  (.D(N_4702_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[45]_net_1 ));
    CFG4 #( .INIT(16'h0906) )  un1_Syn_reg_67_1_a6_2_1 (.A(
        \Parity[0]_net_1 ), .B(\Syn_reg[0]_net_1 ), .C(N_376), .D(
        \un1_Syn_reg[4] ), .Y(un1_Syn_reg_67_1_a6_2_1_net_1));
    CFG4 #( .INIT(16'h8000) )  \Shift_reg_RNI69AG1[2]  (.A(
        \Shift_reg[0]_net_1 ), .B(\Shift_reg[2]_net_1 ), .C(
        \Parity[5]_net_1 ), .D(\Parity[3]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_34));
    CFG4 #( .INIT(16'hB931) )  DataO_6_53_bm (.A(\un22_DataO_i[1] ), 
        .B(DataO_6_53_bm_1_1_net_1), .C(\Shift_reg[24]_net_1 ), .D(
        \Shift_reg[28]_net_1 ), .Y(DataO_6_53_bm_net_1));
    CFG2 #( .INIT(4'h8) )  Shift_reg_1_sqmuxa_1_i_o3_0_a3_1 (.A(
        un14lto4), .B(\Bit_Counter[3]_net_1 ), .Y(N_436_1));
    SLE \TC_Error_Counter[25]  (.D(\TC_Error_Counter_s[25] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[25]));
    SLE \TC_Packet_Counter[9]  (.D(\TC_Packet_Counter_s[9] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[9]));
    SLE \Shift_reg[4]  (.D(N_3580_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[4]_net_1 ));
    SLE \TC_Packet_Counter[11]  (.D(\TC_Packet_Counter_s[11] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[11]));
    CFG4 #( .INIT(16'hB380) )  \un1_block_counter_4[0]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(TC_Packet_Counter18_i_0)
        , .D(un1_block_counter_net_1), .Y(
        \un1_block_counter_4[0]_net_1 ));
    CFG4 #( .INIT(16'h4445) )  Shift_reg_68_37_1293_i_0_2 (.A(
        Shift_reg_68_sn_N_84_mux), .B(
        Shift_reg_68_37_1293_i_0_a2_2_1_net_1), .C(
        \Shift_reg[21]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_37_1293_i_0_2_net_1));
    CFG4 #( .INIT(16'hF780) )  \Shift_reg_68_28[48]  (.A(
        Shift_reg_68_28_6_4), .B(Shift_reg_68_28_3_4), .C(RX_GPIO0_c), 
        .D(\Shift_reg[48]_net_1 ), .Y(N_118));
    CFG4 #( .INIT(16'h195D) )  DataO_10_iv_0_0_RNO_18 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[11]_net_1 ), .D(\Shift_reg[15]_net_1 ), .Y(
        DataO_6_34_1_2));
    CFG4 #( .INIT(16'hC808) )  Shift_reg_68_13_1953_i_i_1_tz (.A(
        N_53_i), .B(\Shift_reg[28]_net_1 ), .C(N_82), .D(N_90), .Y(
        Shift_reg_68_13_1953_i_i_1_tz_net_1));
    CFG4 #( .INIT(16'h503F) )  DataO_10_iv_0_a3_0_RNO_3 (.A(
        \Start_Buff[0]_net_1 ), .B(\Start_Buff[4]_net_1 ), .C(
        \un6_DataO_i[3] ), .D(\un6_DataO_i[2] ), .Y(DataO_2_13_1_2));
    CFG2 #( .INIT(4'h2) )  Shift_reg_68_28_43_0 (.A(N_21_i), .B(N_265), 
        .Y(Shift_reg_68_28_43_0_net_1));
    SLE \TC_Error_Counter[18]  (.D(\TC_Error_Counter_s[18] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[18]));
    CFG4 #( .INIT(16'h78F0) )  Shift_reg_68_61_754_i_m4_am (.A(
        \Shift_reg_68_54_e_0[10] ), .B(Shift_reg_68_54_4), .C(
        \Shift_reg[10]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_61_754_i_m4_am_net_1));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_55_925_i_m4_ns (.A(
        Shift_reg_68_55_925_i_m4_am_net_1), .B(
        Shift_reg_68_55_925_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3583));
    CFG4 #( .INIT(16'h0FAC) )  DataO_10_iv_0_0_RNO_16 (.A(
        \Shift_reg[54]_net_1 ), .B(\Shift_reg[50]_net_1 ), .C(
        DataO_6_10_i_m2_1_2), .D(\Shift_Bit_Counter[5]_net_1 ), .Y(
        N_330));
    CFG2 #( .INIT(4'h8) )  Shift_reg_68_28_9_0 (.A(Shift_reg_68_28_6_4)
        , .B(Shift_reg_68_28_9_2), .Y(Shift_reg_68_28_9_0_net_1));
    CFG3 #( .INIT(8'hD8) )  \Shift_reg_68_28[15]  (.A(
        Shift_reg_68_28_27_net_1), .B(RX_GPIO0_c), .C(
        \Shift_reg[15]_net_1 ), .Y(N_85));
    CFG4 #( .INIT(16'h5410) )  Shift_reg_68_sn_m23_0_a2_RNIC6251 (.A(
        \un1_Syn_reg[0] ), .B(\un1_Syn_reg[6] ), .C(
        Shift_reg_68_sn_N_24), .D(N_53_i), .Y(\Shift_reg_68_54_e_0[8] )
        );
    SLE \Shift_reg[13]  (.D(N_4079_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[13]_net_1 ));
    CFG4 #( .INIT(16'hF0F7) )  un1_State1_1 (.A(N_152), .B(N_356_1), 
        .C(un1_State1_1_0_net_1), .D(TC_Packet_Counter18_i_0), .Y(
        un1_State1_1_net_1));
    CFG4 #( .INIT(16'h0133) )  \un1_block_counter_7_bm[0]  (.A(
        \State1_ns_0_o5_2[0]_net_1 ), .B(Block_ErrO_0_sqmuxa_1_0_net_1)
        , .C(\State1_ns_0_o5_3[0]_net_1 ), .D(
        un1_DataO41_27_a0_0_net_1), .Y(
        \un1_block_counter_7_bm[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[17]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[17]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[16]_net_1 ), .S(
        \TC_Error_Counter_s[17] ), .Y(), .FCO(
        \TC_Error_Counter_cry[17]_net_1 ));
    CFG4 #( .INIT(16'hEFEE) )  Shift_reg_68_6_2159_i_i (.A(N_231), .B(
        N_232), .C(N_217), .D(N_253), .Y(N_59));
    CFG2 #( .INIT(4'h4) )  Shift_reg_68_60_782_i_i_0 (.A(Shift_N_5), 
        .B(Shift_m3_0_a2_2_2), .Y(Shift_reg_68_60_782_i_i_0_net_1));
    CFG3 #( .INIT(8'hF7) )  Shift_reg_68_41_1171_i_o7 (.A(
        \State1[0]_net_1 ), .B(TC_Packet_Counter17_i_0), .C(N_277), .Y(
        N_3793));
    CFG4 #( .INIT(16'h0AFC) )  DataO_10_iv_0_0_RNO_9 (.A(
        \Shift_reg[47]_net_1 ), .B(\Shift_reg[43]_net_1 ), .C(
        \Shift_Bit_Counter[5]_net_1 ), .D(DataO_6_34_1_2), .Y(N_2663));
    SLE \Bit_Counter[4]  (.D(\Bit_Counter_lm[4] ), .CLK(RX_GPIO1_c), 
        .EN(un1_DataO41_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(un14lto4));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIJBE86[16]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[16]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[15] ), .S(
        \TC_Packet_Counter_s[16] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[16] ));
    CFG3 #( .INIT(8'h10) )  \Parity_RNO[5]  (.A(N_2969_1), .B(N_277), 
        .C(N_3723), .Y(N_3720_i_0));
    CFG2 #( .INIT(4'h6) )  \un1_Syn_reg_i_o3[6]  (.A(
        \Syn_reg[6]_net_1 ), .B(\Parity[6]_net_1 ), .Y(
        \un1_Syn_reg[6] ));
    CFG4 #( .INIT(16'h55D5) )  Syn_reg_0_sqmuxa_0 (.A(
        \State1[0]_net_1 ), .B(TC_Packet_Counter17_i_0), .C(N_58), .D(
        N_277), .Y(Syn_reg_0_sqmuxa_0_net_1));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[46]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4680), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4677_i_0));
    CFG4 #( .INIT(16'h8000) )  Shift_reg_68_41_1171_i_a7_0_1 (.A(
        \un1_Syn_reg[0] ), .B(\Shift_reg[25]_net_1 ), .C(N_3793), .D(
        Shift_reg_68_sn_N_82_mux), .Y(
        Shift_reg_68_41_1171_i_a7_0_1_net_1));
    CFG3 #( .INIT(8'hE4) )  Shift_reg_68_36_1321_i_m4 (.A(
        Shift_reg_68_sn_N_84_mux), .B(N_1433_mux), .C(N_1429_mux), .Y(
        N_3913));
    SLE \TC_Error_Counter[0]  (.D(\TC_Error_Counter_s[0] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[0]));
    CFG4 #( .INIT(16'h2112) )  \Syn_reg_RNO[6]  (.A(\Syn_reg[6]_net_1 )
        , .B(N_54), .C(RX_GPIO0_c), .D(\Syn_reg[5]_net_1 ), .Y(
        N_3245_i_0));
    CFG4 #( .INIT(16'h9990) )  \Syn_reg_RNIG6B21[5]  (.A(
        \Syn_reg[5]_net_1 ), .B(\Parity[5]_net_1 ), .C(
        \un1_Syn_reg[3]_net_1 ), .D(\un1_Syn_reg[2] ), .Y(
        Shift_reg_68_sn_N_50));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_10_303_a2 (.A(CCA_NIRQ_c), 
        .B(\Start_Buff[7]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3052));
    CFG3 #( .INIT(8'hFD) )  Shift_reg_68_21_1723_i_i_o2 (.A(
        \Bit_Counter[1]_net_1 ), .B(\Bit_Counter[3]_net_1 ), .C(
        un14lto5), .Y(N_100));
    SLE \TC_Error_Counter[17]  (.D(\TC_Error_Counter_s[17] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[17]));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIONQB5[11]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[11]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[10] ), .S(
        \TC_Packet_Counter_s[11] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[11] ));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_5_358_a2 (.A(CCA_NIRQ_c), .B(
        \Start_Buff[2]_net_1 ), .C(\State1[0]_net_1 ), .Y(
        Start_Buff_10_5_358_a2_net_1));
    CFG2 #( .INIT(4'h8) )  un1_DataO41_22_0_a3_0_3 (.A(N_298), .B(
        N_94_i), .Y(un1_DataO41_22_0_a3_0_2));
    CFG4 #( .INIT(16'hEFE0) )  Shift_reg_68_1_2300_i_0_m3 (.A(N_86), 
        .B(Shift_reg_68_1_2300_i_0_o3_1_0_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .D(N_392), .Y(N_403));
    CFG3 #( .INIT(8'h40) )  Shift_reg_68_19_1783_i_0_a2_2_1_0 (.A(
        N_381), .B(\Shift_reg[34]_net_1 ), .C(N_417_1), .Y(
        Shift_reg_68_19_1783_i_0_a2_2_1_net_1));
    CFG4 #( .INIT(16'h4000) )  \Shift_reg_RNO_2[43]  (.A(
        \un1_Syn_reg[2] ), .B(N_53_i), .C(\un1_Syn_reg[0] ), .D(
        \un1_Syn_reg[6] ), .Y(\Shift_reg_RNO_2[43]_net_1 ));
    CFG4 #( .INIT(16'h0545) )  Start_Buff_0_sqmuxa_0_0_RNIEMTP1 (.A(
        un1_CCA_i_0), .B(N_277), .C(Start_Buff_0_sqmuxa_0_0_net_1), .D(
        un1_DataO41_26_i_1), .Y(un1_DataO41_26_i_0));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_6_347_a2 (.A(CCA_NIRQ_c), .B(
        \Start_Buff[3]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3092));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIB04N3[6]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[6]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Packet_Counter_cry[5] ), .S(
        \TC_Packet_Counter_s[6] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[6] ));
    SLE \Bit_Counter[5]  (.D(\Bit_Counter_lm[5] ), .CLK(RX_GPIO1_c), 
        .EN(un1_DataO41_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(un14lto5));
    CFG4 #( .INIT(16'h0004) )  \Shift_reg_RNIR9GB1[55]  (.A(
        \Parity[1]_net_1 ), .B(\Shift_reg[55]_net_1 ), .C(
        \Parity[6]_net_1 ), .D(\Parity[0]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_32));
    CFG3 #( .INIT(8'h7F) )  DataO_10_iv_0_o2 (.A(
        \Shift_Bit_Counter[3]_net_1 ), .B(\Shift_Bit_Counter[5]_net_1 )
        , .C(\Shift_Bit_Counter[4]_net_1 ), .Y(N_302));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[1]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3655), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3652_i_0));
    CFG4 #( .INIT(16'h1131) )  Shift_reg_68_29_1522_i_a7 (.A(
        \State1[0]_net_1 ), .B(\Shift_reg[13]_net_1 ), .C(
        Shift_reg_68_sn_N_73), .D(un1_TC_Packet_Counter17_3_net_1), .Y(
        N_4080));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_35_1349_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_82), 
        .D(N_89), .Y(N_3940));
    SLE \Shift_reg[51]  (.D(N_4558_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[51]_net_1 ));
    CFG4 #( .INIT(16'h0B00) )  \Shift_reg_RNO[13]  (.A(N_1451_mux), .B(
        N_349_1), .C(N_4084), .D(N_4079_i_1), .Y(N_4079_i_0));
    CFG4 #( .INIT(16'hF0E2) )  Parity_16_0_1066_i_m5 (.A(RX_GPIO0_c), 
        .B(\Parity_Counter[0]_net_1 ), .C(\Parity[6]_net_1 ), .D(
        N_3721), .Y(N_3703));
    CFG4 #( .INIT(16'h9009) )  \Syn_reg_RNIUMFH1_1[3]  (.A(
        \Syn_reg[3]_net_1 ), .B(\Parity[3]_net_1 ), .C(
        \Syn_reg[2]_net_1 ), .D(\Parity[2]_net_1 ), .Y(
        Shift_reg_68_sn_N_9));
    CFG4 #( .INIT(16'h1000) )  \State1_ns_0_a5_1[0]  (.A(
        \block_counter[0]_net_1 ), .B(\block_counter[1]_net_1 ), .C(
        \State1_ns_0_a5_1_0[0]_net_1 ), .D(\State1[0]_net_1 ), .Y(
        N_2130));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[24]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3819), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3816_i_0));
    CFG4 #( .INIT(16'hE323) )  DataO_10_iv_0_0_RNO_6 (.A(N_1074), .B(
        DataO_6_15_1_2), .C(\un22_DataO_i[0] ), .D(N_330), .Y(N_2644));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_1_657_a2 (.A(CCA_NIRQ_c), .B(
        \Start_Buff[14]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3346));
    CFG2 #( .INIT(4'h4) )  un1_DataO41_27_a0_0 (.A(un1_DataI), .B(
        TC_Packet_Counter17_i_0), .Y(un1_DataO41_27_a0_0_net_1));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_4_2216_i_m4_ns (.A(
        Shift_reg_68_4_2216_i_m4_am_net_1), .B(
        Shift_reg_68_4_2216_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4655));
    CFG4 #( .INIT(16'hC400) )  Shift_reg_68_30_1493_i_i_o3_1_0_RNO (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(TC_Packet_Counter17_i_0)
        , .D(N_102), .Y(Shift_m5_0));
    CFG3 #( .INIT(8'h12) )  \Parity_Counter_9[1]  (.A(CO0_0), .B(
        \un1_block_counter_4[0]_net_1 ), .C(\Parity_Counter[1]_net_1 ), 
        .Y(\Parity_Counter_9[1]_net_1 ));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_17_1839_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(N_82), .C(Shift_reg_68_sn_N_84_mux), 
        .D(N_102_0), .Y(N_4347));
    SLE \Shift_reg[27]  (.D(N_69), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[27]_net_1 ));
    SLE \Shift_reg[43]  (.D(N_4752_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[43]_net_1 ));
    CFG4 #( .INIT(16'h0AFC) )  DataO_10_iv_0_0_RNO_14 (.A(
        \Shift_reg[52]_net_1 ), .B(\Shift_reg[48]_net_1 ), .C(
        \Shift_Bit_Counter[5]_net_1 ), .D(DataO_6_13_i_m2_1_2), .Y(
        N_1074));
    CFG4 #( .INIT(16'h0AFC) )  DataO_10_iv_0_0_RNO_20 (.A(
        \Shift_reg[39]_net_1 ), .B(\Shift_reg[35]_net_1 ), .C(
        \Shift_Bit_Counter[5]_net_1 ), .D(DataO_6_18_i_m2_1_2), .Y(
        N_325));
    SLE \TC_Packet_Counter[15]  (.D(\TC_Packet_Counter_s[15] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[15]));
    CFG4 #( .INIT(16'h0A02) )  State2_1_sqmuxa (.A(CCA_NIRQ_c), .B(
        \State2[0]_net_1 ), .C(\State2[1]_net_1 ), .D(N_302), .Y(
        State2_1_sqmuxa_net_1));
    CFG4 #( .INIT(16'h0B00) )  \Shift_reg_RNO[3]  (.A(N_1426_mux), .B(
        N_349_1), .C(N_3610), .D(N_3605_i_1), .Y(N_3605_i_0));
    ARI1 #( .INIT(20'h4AA00) )  Bit_Counter_s_369 (.A(VCC_net_1), .B(
        un14lto0), .C(GND_net_1), .D(GND_net_1), .FCI(VCC_net_1), .S(), 
        .Y(), .FCO(Bit_Counter_s_369_FCO));
    CFG3 #( .INIT(8'h08) )  un39_Shift_reg_0 (.A(
        \Bit_Counter[1]_net_1 ), .B(\Bit_Counter[2]_net_1 ), .C(
        un14lto0), .Y(un39_Shift_reg_0_net_1));
    SLE \TC_Error_Counter[26]  (.D(\TC_Error_Counter_s[26] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[26]));
    CFG4 #( .INIT(16'h888A) )  Shift_reg_68_6_2159_i_i_a2_3 (.A(
        Shift_reg_68_6_2159_i_i_a2_3_2_net_1), .B(
        un1_TC_Packet_Counter17_3_net_1), .C(Shift_N_7_1), .D(
        Shift_reg_68_sn_N_73), .Y(N_253));
    SLE \TC_Error_Counter[21]  (.D(\TC_Error_Counter_s[21] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[21]));
    CFG3 #( .INIT(8'h1B) )  Shift_reg_68_37_1293_i_0_1_1 (.A(N_402), 
        .B(RX_GPIO0_c), .C(\Shift_reg[21]_net_1 ), .Y(
        Shift_reg_68_37_1293_i_0_1_1_net_1));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[55]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4467), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4464_i_0));
    SLE \Shift_reg[5]  (.D(N_3558_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[5]_net_1 ));
    CFG4 #( .INIT(16'h32FA) )  \Shift_reg_RNO_0[53]  (.A(
        \Shift_reg[53]_net_1 ), .B(\State1[0]_net_1 ), .C(
        Shift_reg_68_sn_N_84_mux), .D(un1_TC_Packet_Counter17_5_net_1), 
        .Y(N_4511_i_1));
    CFG3 #( .INIT(8'h5D) )  Shift_reg_68_1_2300_i_0_o2_0 (.A(
        CCA_NIRQ_c), .B(\State1[0]_net_1 ), .C(TC_Packet_Counter17_i_0)
        , .Y(Shift_reg_68_1_2300_i_0_o2));
    ARI1 #( .INIT(20'h4A200) )  un1_DataO41_18_1_0_RNIGFRM (.A(
        VCC_net_1), .B(N_3002), .C(TC_Packet_Counter17_i_0), .D(N_277), 
        .FCI(VCC_net_1), .S(), .Y(un1_DataO41_18_1_0_RNIGFRM_Y), .FCO(
        TC_Packet_Counter_cry_cy));
    CFG4 #( .INIT(16'hFB40) )  Shift_reg_68_59_810_i_m4_bm (.A(N_34), 
        .B(Shift_reg_68_28_3_4), .C(RX_GPIO0_c), .D(
        \Shift_reg[8]_net_1 ), .Y(Shift_reg_68_59_810_i_m4_bm_net_1));
    CFG3 #( .INIT(8'hFE) )  un1_Syn_reg_2_0_a3_RNINA0E1 (.A(
        un1_Syn_reg_2), .B(N_2847), .C(N_2846), .Y(
        un1_Syn_reg_2_0_a3_RNINA0E1_net_1));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_14_259_a2 (.A(CCA_NIRQ_c), 
        .B(\Start_Buff[11]_net_1 ), .C(\State1[0]_net_1 ), .Y(
        Start_Buff_10_14_259_a2_net_1));
    SLE Enable (.D(\Shift_Bit_Counter_cry_cy_Y[0] ), .CLK(RX_GPIO1_c), 
        .EN(un1_DataO41_8_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(ENASM_0));
    CFG4 #( .INIT(16'hF780) )  Shift_reg_68_27_1552_i_m4_bm (.A(
        Shift_reg_68_28_25_4), .B(Shift_reg_68_28_50_4), .C(RX_GPIO0_c)
        , .D(\Shift_reg[42]_net_1 ), .Y(
        Shift_reg_68_27_1552_i_m4_bm_net_1));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[19]  (.A(
        Shift_reg_68_28_31_0_net_1), .B(N_92), .C(RX_GPIO0_c), .D(
        \Shift_reg[19]_net_1 ), .Y(N_89));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[24]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[24]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[23]_net_1 ), .S(
        \TC_Error_Counter_s[24] ), .Y(), .FCO(
        \TC_Error_Counter_cry[24]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \Shift_Bit_Counter_s[5]  (.A(VCC_net_1)
        , .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_Bit_Counter_cry_cy_Y[0] ), .D(GND_net_1), .FCI(
        \Shift_Bit_Counter_cry[4]_net_1 ), .S(
        \Shift_Bit_Counter_s[5]_net_1 ), .Y(), .FCO());
    CFG2 #( .INIT(4'h7) )  un1_TC_Packet_Counter17_1 (.A(N_277), .B(
        TC_Packet_Counter17_i_0), .Y(un1_TC_Packet_Counter17_1_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[3]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[3]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[2]_net_1 ), .S(
        \TC_Error_Counter_s[3] ), .Y(), .FCO(
        \TC_Error_Counter_cry[3]_net_1 ));
    CFG4 #( .INIT(16'h0008) )  un1_Start_Buff_1_6 (.A(
        \Start_Buff[8]_net_1 ), .B(\Start_Buff[7]_net_1 ), .C(
        \Start_Buff[6]_net_1 ), .D(\Start_Buff[5]_net_1 ), .Y(
        un1_Start_Buff_1_6_net_1));
    CFG3 #( .INIT(8'h02) )  Shift_reg_68_28_8_0 (.A(
        Shift_reg_68_28_6_4), .B(\Bit_Counter[2]_net_1 ), .C(un14lto0), 
        .Y(Shift_reg_68_28_8_0_net_1));
    CFG2 #( .INIT(4'hD) )  Shift_reg_68_28_20_1_o3 (.A(un14lto4), .B(
        \Bit_Counter[1]_net_1 ), .Y(N_110));
    ARI1 #( .INIT(20'h48800) )  \Shift_Bit_Counter_cry[3]  (.A(
        VCC_net_1), .B(\Shift_Bit_Counter[3]_net_1 ), .C(
        \Shift_Bit_Counter_cry_cy_Y[0] ), .D(GND_net_1), .FCI(
        \Shift_Bit_Counter_cry[2]_net_1 ), .S(\Shift_Bit_Counter_s[3] )
        , .Y(), .FCO(\Shift_Bit_Counter_cry[3]_net_1 ));
    CFG4 #( .INIT(16'hAAA8) )  Shift_reg_68_63_697_i_i_a2_0_1 (.A(
        \Shift_reg[12]_net_1 ), .B(\Bit_Counter[2]_net_1 ), .C(N_103), 
        .D(N_86), .Y(Shift_reg_68_63_697_i_i_a2_0));
    CFG3 #( .INIT(8'h10) )  \Parity_RNO[0]  (.A(N_2969_1), .B(N_277), 
        .C(N_275), .Y(N_3227_i_0));
    SLE \Bit_Counter[0]  (.D(\Bit_Counter_lm[0] ), .CLK(RX_GPIO1_c), 
        .EN(un1_DataO41_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(un14lto0));
    SLE \TC_Packet_Counter[31]  (.D(\TC_Packet_Counter_s[31] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[31]));
    CFG4 #( .INIT(16'hF8FF) )  Shift_reg_68_28_12_1_i_o2 (.A(N_436_1), 
        .B(un14lto5), .C(Shift_reg_68_28_12_1_i_o2_1_net_1), .D(
        TC_Packet_Counter17_i_0), .Y(N_86));
    CFG4 #( .INIT(16'hFF80) )  DataO_10_iv_0_0 (.A(N_302), .B(
        DataO_10_iv_0_a3_0_net_1), .C(N_309), .D(N_354), .Y(DataO_10));
    CFG4 #( .INIT(16'h3337) )  Shift_reg_68_29_1522_i_0 (.A(
        \Shift_reg[13]_net_1 ), .B(CCA_NIRQ_c), .C(
        Shift_reg_68_sn_N_56), .D(N_82), .Y(
        Shift_reg_68_29_1522_i_0_net_1));
    SLE \TC_Packet_Counter[27]  (.D(\TC_Packet_Counter_s[27] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[27]));
    CFG4 #( .INIT(16'h3337) )  Shift_reg_68_11_2010_i_0 (.A(
        \Shift_reg[54]_net_1 ), .B(CCA_NIRQ_c), .C(
        Shift_reg_68_sn_N_56), .D(N_82), .Y(
        Shift_reg_68_11_2010_i_0_net_1));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_61_754_i_m4_ns (.A(
        Shift_reg_68_61_754_i_m4_am_net_1), .B(
        Shift_reg_68_61_754_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3436));
    CFG4 #( .INIT(16'h5030) )  \un1_Syn_reg_i_o3_0_x2_RNI64E57[1]  (.A(
        Shift_reg_68_sn_m59_i_x3_RNI3Q7P3_net_1), .B(
        Shift_reg_68_sn_m72_6_ns_1), .C(N_53_i), .D(\un1_Syn_reg[6] ), 
        .Y(Shift_reg_68_sn_m72_7_ns_sx));
    CFG4 #( .INIT(16'h0010) )  \Shift_reg_RNO[22]  (.A(N_3868), .B(
        N_3863_i_1_1), .C(N_3863_i_1), .D(N_3866), .Y(N_3863_i_0));
    CFG4 #( .INIT(16'h2303) )  IP_END_RNO (.A(\State1[0]_net_1 ), .B(
        un1_CCA_i_0), .C(Start_Buff_0_sqmuxa_1_net_1), .D(
        TC_Packet_Counter19_net_1), .Y(un1_DataO41_19_i_0));
    CFG4 #( .INIT(16'h0F53) )  DataO_6_53_bm_1_1 (.A(
        \Shift_reg[26]_net_1 ), .B(\Shift_reg[30]_net_1 ), .C(
        \un22_DataO_i[2] ), .D(\un22_DataO_i[1] ), .Y(
        DataO_6_53_bm_1_1_net_1));
    CFG4 #( .INIT(16'h0007) )  \Shift_reg_RNO[50]  (.A(
        \State1[0]_net_1 ), .B(un1_TC_Packet_Counter17_5_net_1), .C(
        N_4585), .D(Shift_reg_68_7_2129_i_2_net_1), .Y(N_4580_i_0));
    CFG3 #( .INIT(8'hD8) )  Shift_reg_68_47_1039_i_m4_0_ns (.A(N_82), 
        .B(Shift_reg_68_47_1039_i_m4_0_bm_net_1), .C(
        Shift_reg_68_47_1039_i_m4_0_am_net_1), .Y(N_3679));
    SLE \Shift_reg[21]  (.D(N_3885_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[21]_net_1 ));
    SLE \Shift_Bit_Counter[0]  (.D(\Shift_Bit_Counter_s[0] ), .CLK(
        RX_GPIO1_c), .EN(Shift_Bit_Countere), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \un22_DataO_i[0] ));
    CFG3 #( .INIT(8'h04) )  \Shift_reg_RNO[19]  (.A(
        Shift_reg_68_35_1349_i_1_net_1), .B(N_3935_i_1), .C(N_3940), 
        .Y(N_3935_i_0));
    CFG2 #( .INIT(4'hB) )  un1_DataO41_8_0_o2 (.A(
        TC_Packet_Counter17_i_0), .B(\State1[0]_net_1 ), .Y(N_305));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNISM365[10]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[10]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[9] ), .S(
        \TC_Packet_Counter_s[10] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[10] ));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[0]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3680), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3677_i_0));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_56_895_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_82), 
        .D(N_75_0), .Y(N_3563));
    SLE \Syn_reg[6]  (.D(N_3245_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_15_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Syn_reg[6]_net_1 ));
    CFG4 #( .INIT(16'h00C4) )  Shift_reg_68_13_1953_i_i_o3_0 (.A(
        N_94_i), .B(Shift_reg_68_13_1953_i_i_o3_0_0_0), .C(N_82), .D(
        Shift_N_7_mux_2), .Y(Shift_reg_68_13_1953_i_i_o3_0_0_net_1));
    SLE \TC_Error_Counter[19]  (.D(\TC_Error_Counter_s[19] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[19]));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_32_1435_i_m4_ns (.A(
        Shift_reg_68_32_1435_i_m4_am_net_1), .B(
        Shift_reg_68_32_1435_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4010));
    CFG4 #( .INIT(16'hFFFE) )  un1_Syn_reg_2_0_a3_RNIEDI03 (.A(
        un1_Syn_reg_2), .B(N_2847), .C(N_2846), .D(N_2843), .Y(
        Shift_m4_e_1_sx));
    SLE \Shift_reg[17]  (.D(N_3982_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[17]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIS3KP6[19]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[19]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[18] ), .S(
        \TC_Packet_Counter_s[19] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[19] ));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[35]  (.A(
        Shift_reg_68_28_17_0_net_1), .B(N_92), .C(RX_GPIO0_c), .D(
        \Shift_reg[35]_net_1 ), .Y(N_105));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_40_1205_i_m4_ns (.A(
        Shift_reg_68_40_1205_i_m4_am_net_1), .B(
        Shift_reg_68_40_1205_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3819));
    SLE \State1[0]  (.D(\State1_ns[0] ), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\State1[0]_net_1 ));
    CFG4 #( .INIT(16'h6A00) )  Shift_reg_68_21_1723_i_i_a2_2_0 (.A(
        \Shift_reg[36]_net_1 ), .B(Shift_reg_68_43_2), .C(
        Shift_reg_68_50_net_1), .D(Shift_reg_68_sn_N_56), .Y(
        Shift_reg_68_21_1723_i_i_a2_2_0_net_1));
    CFG4 #( .INIT(16'h4000) )  Shift_reg_68_28_30_0 (.A(un14lto4), .B(
        \Bit_Counter[2]_net_1 ), .C(un14lto5), .D(Shift_reg_68_28_30_3)
        , .Y(Shift_reg_68_28_30_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[15]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[15]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[14]_net_1 ), .S(
        \TC_Error_Counter_s[15] ), .Y(), .FCO(
        \TC_Error_Counter_cry[15]_net_1 ));
    SLE \Parity[1]  (.D(N_3207_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_10_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Parity[1]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \Shift_reg_RNIISG6[24]  (.A(
        \Shift_reg[30]_net_1 ), .B(\Shift_reg[24]_net_1 ), .C(
        \Shift_reg[23]_net_1 ), .D(\Shift_reg[22]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_37));
    CFG2 #( .INIT(4'h6) )  \un1_Syn_reg[3]  (.A(\Parity[3]_net_1 ), .B(
        \Syn_reg[3]_net_1 ), .Y(\un1_Syn_reg[3]_net_1 ));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[11]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3411), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3408_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[19]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[19]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[18]_net_1 ), .S(
        \TC_Error_Counter_s[19] ), .Y(), .FCO(
        \TC_Error_Counter_cry[19]_net_1 ));
    CFG3 #( .INIT(8'h8A) )  Syn_reg_0_sqmuxa_2 (.A(CCA_NIRQ_c), .B(
        \State1[0]_net_1 ), .C(un1_Start_Buff_1_net_1), .Y(
        Syn_reg_0_sqmuxa_2_net_1));
    CFG4 #( .INIT(16'h0001) )  \Shift_reg_RNIP4I6[20]  (.A(
        \Shift_reg[29]_net_1 ), .B(\Shift_reg[45]_net_1 ), .C(
        \Shift_reg[21]_net_1 ), .D(\Shift_reg[20]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_46));
    SLE \Syn_reg[1]  (.D(N_3319_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_15_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Syn_reg[1]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \State1_ns_0_o5[0]  (.A(
        \State1_ns_0_o5_3[0]_net_1 ), .B(\State1_ns_0_o5_2[0]_net_1 ), 
        .Y(N_2121));
    CFG4 #( .INIT(16'hB931) )  DataO_10_iv_0_a3_0_RNO_1 (.A(
        \un6_DataO_i[2] ), .B(DataO_2_10_1_2), .C(
        \Start_Buff[2]_net_1 ), .D(\Start_Buff[10]_net_1 ), .Y(N_2624));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIHG302[2]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[2]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Packet_Counter_cry[1] ), .S(
        \TC_Packet_Counter_s[2] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[2] ));
    SLE \Shift_Bit_Counter[1]  (.D(\Shift_Bit_Counter_s[1] ), .CLK(
        RX_GPIO1_c), .EN(Shift_Bit_Countere), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \un22_DataO_i[1] ));
    CFG2 #( .INIT(4'hB) )  Shift_reg_68_60_782_i_i_o2_0 (.A(N_91), .B(
        un14lto5), .Y(N_103));
    CFG4 #( .INIT(16'h840C) )  Shift_reg_68_7_2129_i_a7_1_0 (.A(
        Shift_reg_68_50_2), .B(Shift_reg_68_sn_N_56), .C(
        \Shift_reg[50]_net_1 ), .D(\un1_Syn_reg[0] ), .Y(
        Shift_reg_68_7_2129_i_a7_1_0_net_1));
    CFG4 #( .INIT(16'h0001) )  \Shift_reg_RNIISKN[11]  (.A(
        \Shift_reg[17]_net_1 ), .B(\Shift_reg[11]_net_1 ), .C(
        \Shift_reg[5]_net_1 ), .D(\Shift_reg[3]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_42));
    CFG4 #( .INIT(16'hF078) )  Shift_reg_68_25_1609_i_m4_am (.A(
        \Shift_reg_68_54_e_0[10] ), .B(Shift_reg_68_54_4), .C(
        \Shift_reg[40]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_25_1609_i_m4_am_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[30]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[30]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[29]_net_1 ), .S(
        \TC_Error_Counter_s[30] ), .Y(), .FCO(
        \TC_Error_Counter_cry[30]_net_1 ));
    CFG4 #( .INIT(16'h00B8) )  un1_DataO41_22_0_1 (.A(N_3002), .B(
        un1_DataI), .C(un1_DataO41_22_0_a3_1), .D(
        un1_TC_Packet_Counter17_1_net_1), .Y(un1_DataO41_22_0_1_net_1));
    CFG2 #( .INIT(4'h4) )  \Syn_reg_RNO[5]  (.A(N_54), .B(
        \Syn_reg[4]_net_1 ), .Y(N_3263_i_0));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_13_270_a2 (.A(CCA_NIRQ_c), 
        .B(\Start_Buff[10]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3022));
    CFG2 #( .INIT(4'hD) )  Shift_reg_68_30_1493_i_i_o2 (.A(un14lto5), 
        .B(\Bit_Counter[1]_net_1 ), .Y(N_102));
    SLE \TC_Packet_Counter[1]  (.D(\TC_Packet_Counter_s[1] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[1]));
    CFG3 #( .INIT(8'hD8) )  Shift_reg_68_16_1869_i_m4_bm (.A(
        Shift_reg_68_28_13_net_1), .B(RX_GPIO0_c), .C(
        \Shift_reg[31]_net_1 ), .Y(Shift_reg_68_16_1869_i_m4_bm_net_1));
    SLE \TC_Packet_Counter[19]  (.D(\TC_Packet_Counter_s[19] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[19]));
    SLE \Shift_reg[11]  (.D(N_3408_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[11]_net_1 ));
    CFG4 #( .INIT(16'h0310) )  Shift_reg_68_50 (.A(\un1_Syn_reg[2] ), 
        .B(N_53_i), .C(\un1_Syn_reg[0] ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_50_net_1));
    CFG4 #( .INIT(16'h195D) )  DataO_10_iv_0_0_RNO_28 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[1]_net_1 ), .D(\Shift_reg[5]_net_1 ), .Y(
        DataO_6_21_i_m2_1_2));
    CFG3 #( .INIT(8'h10) )  \Parity_RNO[1]  (.A(N_2969_1), .B(N_277), 
        .C(N_80), .Y(N_3207_i_0));
    CFG4 #( .INIT(16'h5030) )  \un1_Syn_reg_i_o3_0_x2_RNI64E57_0[1]  (
        .A(Shift_reg_68_sn_m59_i_x3_RNI3Q7P3_net_1), .B(
        Shift_reg_68_sn_m72_6_ns_1), .C(N_53_i), .D(\un1_Syn_reg[6] ), 
        .Y(Shift_m3_0_sx_sx));
    SLE \Start_Buff[9]  (.D(N_3042), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[9]_net_1 ));
    CFG4 #( .INIT(16'hFF40) )  \State1_ns_0[0]  (.A(
        un1_TC_Packet_Counter17_3_net_1), .B(N_3002), .C(N_2121), .D(
        \State1_ns_0_1[0]_net_1 ), .Y(\State1_ns[0] ));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[3]  (.A(
        Shift_reg_68_28_43_0_net_1), .B(N_92), .C(RX_GPIO0_c), .D(
        \Shift_reg[3]_net_1 ), .Y(N_73_0));
    SLE \Shift_reg[47]  (.D(N_4652_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[47]_net_1 ));
    CFG3 #( .INIT(8'hF7) )  Shift_reg_68_28_0_i_0 (.A(
        \Bit_Counter[1]_net_1 ), .B(\State1[0]_net_1 ), .C(N_58), .Y(
        N_374));
    CFG4 #( .INIT(16'h8880) )  un1_DataO41_22_0_a3_1_0 (.A(N_3002), .B(
        N_244_2), .C(N_373), .D(N_372), .Y(un1_DataO41_22_0_a3_1));
    CFG4 #( .INIT(16'hF600) )  \Syn_reg_RNIPJ811[1]  (.A(
        \Parity[1]_net_1 ), .B(\Syn_reg[1]_net_1 ), .C(
        \un1_Syn_reg[5] ), .D(\State1[0]_net_1 ), .Y(
        Shift_reg_68_sn_N_78_mux));
    CFG4 #( .INIT(16'hFA3A) )  Shift_reg_68_sn_m21_0_a2_0_x2_RNIV2771 
        (.A(N_97_i), .B(\un1_Syn_reg[3]_net_1 ), .C(\un1_Syn_reg[0] ), 
        .D(\un1_Syn_reg[2] ), .Y(Shift_reg_68_sn_N_32));
    SLE \TC_Error_Counter[30]  (.D(\TC_Error_Counter_s[30] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[30]));
    CFG4 #( .INIT(16'h0660) )  un1_Syn_reg_2_0_a2_0 (.A(
        \Parity[5]_net_1 ), .B(\Syn_reg[5]_net_1 ), .C(
        \Syn_reg[6]_net_1 ), .D(\Parity[6]_net_1 ), .Y(N_94_i));
    CFG2 #( .INIT(4'h2) )  Shift_reg_68_sn_m57_i_o3_RNIB4CN (.A(
        Shift_reg_68_sn_N_16), .B(\un1_Syn_reg[5] ), .Y(
        \Shift_reg_68_54_e_0[4] ));
    CFG4 #( .INIT(16'h195D) )  DataO_10_iv_0_0_RNO_26 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[18]_net_1 ), .D(\Shift_reg[22]_net_1 ), .Y(
        DataO_6_10_i_m2_1_2));
    CFG2 #( .INIT(4'h8) )  \State1_ns_0_a5_2_1[0]  (.A(
        \Start_Buff[4]_net_1 ), .B(CCA_NIRQ_c), .Y(N_2131_1));
    CFG3 #( .INIT(8'hD8) )  \un1_Syn_reg_RNIQLBC[3]  (.A(
        \un1_Syn_reg[2] ), .B(\un1_Syn_reg[5] ), .C(
        \un1_Syn_reg[3]_net_1 ), .Y(\un1_Syn_reg_RNIQLBC[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[5]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[5]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[4]_net_1 ), .S(
        \TC_Error_Counter_s[5] ), .Y(), .FCO(
        \TC_Error_Counter_cry[5]_net_1 ));
    CFG4 #( .INIT(16'hF078) )  Shift_reg_68_42_1143_i_m4_am (.A(
        \Shift_reg_68_54_e_0[26] ), .B(Shift_reg_68_54_net_1), .C(
        \Shift_reg[26]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_42_1143_i_m4_am_net_1));
    CFG4 #( .INIT(16'hF780) )  Shift_reg_68_25_1609_i_m4_bm (.A(
        Shift_reg_68_28_22_1_net_1), .B(Shift_reg_68_28_3_4), .C(
        RX_GPIO0_c), .D(\Shift_reg[40]_net_1 ), .Y(
        Shift_reg_68_25_1609_i_m4_bm_net_1));
    SLE \Syn_reg[0]  (.D(N_3332_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_15_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Syn_reg[0]_net_1 ));
    CFG4 #( .INIT(16'hFFBF) )  un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_sx (.A(
        \Shift_reg[53]_net_1 ), .B(\Parity[4]_net_1 ), .C(
        \Parity[2]_net_1 ), .D(\Shift_reg[51]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_sx_net_1));
    CFG4 #( .INIT(16'h530F) )  DataO_10_iv_0_a3_0_RNO_7 (.A(
        \Start_Buff[1]_net_1 ), .B(\Start_Buff[5]_net_1 ), .C(
        \un6_DataO_i[2] ), .D(\un6_DataO_i[3] ), .Y(DataO_2_6_1_2));
    CFG2 #( .INIT(4'h8) )  un1_DataO41_18_1_0 (.A(\State1[0]_net_1 ), 
        .B(CCA_NIRQ_c), .Y(N_3002));
    CFG4 #( .INIT(16'h0002) )  Shift_reg_68_57_866_i_i_a2_3_1 (.A(
        Shift_reg_68_57_866_i_i_a2_3_1_1_net_1), .B(
        Shift_reg_68_sn_N_56), .C(\Shift_reg[6]_net_1 ), .D(N_123), .Y(
        Shift_reg_68_57_866_i_i_a2_3_1_net_1));
    SLE \Parity_Counter[0]  (.D(\Parity_Counter_9[0]_net_1 ), .CLK(
        RX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Parity_Counter[0]_net_1 ));
    CFG4 #( .INIT(16'h0010) )  \Shift_reg_RNO[53]  (.A(N_4516), .B(
        N_4511_i_1_1), .C(N_4511_i_1), .D(N_4514), .Y(N_4511_i_0));
    SLE \Shift_reg[52]  (.D(N_4533_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[52]_net_1 ));
    CFG4 #( .INIT(16'h0660) )  un1_Syn_reg_2_0_a2 (.A(
        \Syn_reg[4]_net_1 ), .B(\Parity[4]_net_1 ), .C(
        \Syn_reg[2]_net_1 ), .D(\Parity[2]_net_1 ), .Y(N_370));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[4]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[4]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[3]_net_1 ), .S(
        \TC_Error_Counter_s[4] ), .Y(), .FCO(
        \TC_Error_Counter_cry[4]_net_1 ));
    CFG3 #( .INIT(8'h08) )  DataO_10_iv_0_a3_0 (.A(DataO_2), .B(
        DataO_0_sqmuxa_1_0_net_1), .C(TC_Packet_Counter18_i_0), .Y(
        N_354));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_51_1011_i_m4_ns (.A(
        Shift_reg_68_51_1011_i_m4_am_net_1), .B(
        Shift_reg_68_51_1011_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3655));
    CFG3 #( .INIT(8'hD8) )  Shift_reg_68_40_1205_i_m4_bm (.A(
        Shift_reg_68_28_36_net_1), .B(RX_GPIO0_c), .C(
        \Shift_reg[24]_net_1 ), .Y(Shift_reg_68_40_1205_i_m4_bm_net_1));
    CFG3 #( .INIT(8'hF7) )  Shift_reg_68_46_1115_i_i_N_7L14 (.A(
        Shift_reg_68_54_4), .B(Shift_reg_68_46_1115_i_i_N_4L7_net_1), 
        .C(\un1_Syn_reg[0] ), .Y(Shift_reg_68_46_1115_i_i_N_7L14_net_1)
        );
    SLE \TC_Error_Counter[22]  (.D(\TC_Error_Counter_s[22] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[22]));
    CFG3 #( .INIT(8'h13) )  Shift_reg_68_41_1171_i_a7_0_0 (.A(
        Shift_reg_68_sn_N_82_mux), .B(\Shift_reg[25]_net_1 ), .C(
        \un1_Syn_reg[0] ), .Y(Shift_reg_68_41_1171_i_a7_0));
    CFG3 #( .INIT(8'hE2) )  DataO_6_53_ns (.A(DataO_6_53_am_net_1), .B(
        \un22_DataO_i[0] ), .C(DataO_6_53_bm_net_1), .Y(N_2682));
    CFG4 #( .INIT(16'h3337) )  Shift_reg_68_39_1233_i_0 (.A(
        \Shift_reg[23]_net_1 ), .B(CCA_NIRQ_c), .C(
        Shift_reg_68_sn_N_56), .D(N_82), .Y(
        Shift_reg_68_39_1233_i_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIJCSA7[22]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[22]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[21] ), .S(
        \TC_Packet_Counter_s[22] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[22] ));
    CFG2 #( .INIT(4'h2) )  Shift_reg_68_28_15_1 (.A(
        Shift_reg_68_28_29_3), .B(un14lto5), .Y(
        Shift_reg_68_28_15_0_net_1));
    CFG4 #( .INIT(16'h1110) )  un1_TC_Packet_Counter17_3_RNI29NGA (.A(
        Shift_m3_0_sx_sx), .B(un1_TC_Packet_Counter17_3_net_1), .C(
        N_53_i), .D(N_2548), .Y(Shift_m3_0_sx));
    CFG3 #( .INIT(8'h9A) )  Shift_reg_68_62_726_i_m4_am (.A(
        \Shift_reg[11]_net_1 ), .B(\un1_Syn_reg[6] ), .C(N_1435), .Y(
        Shift_reg_68_62_726_i_m4_am_net_1));
    CFG4 #( .INIT(16'h0800) )  \Parity_Counter_RNI1GJT[0]  (.A(
        \Parity_Counter[0]_net_1 ), .B(\State1[0]_net_1 ), .C(
        un1_CCA_i_0), .D(N_58), .Y(CO0_0));
    CFG2 #( .INIT(4'hE) )  un1_DataO41_22_0_o2 (.A(\un1_Syn_reg[0] ), 
        .B(N_53_i), .Y(N_298));
    CFG2 #( .INIT(4'h8) )  \Bit_Counter_lm_0[2]  (.A(
        Bit_Counter_3_sqmuxa), .B(\Bit_Counter_s[2] ), .Y(
        \Bit_Counter_lm[2] ));
    CFG4 #( .INIT(16'h6996) )  un1_Syn_reg_67_1_x2_1_a3_0_x3 (.A(
        \un1_Syn_reg[2] ), .B(\un1_Syn_reg[3]_net_1 ), .C(
        \un1_Syn_reg[6] ), .D(\un1_Syn_reg[5] ), .Y(N_73_i));
    CFG3 #( .INIT(8'hFE) )  Shift_reg_68_28_0_a3_0_o3 (.A(
        \Bit_Counter[2]_net_1 ), .B(un14lto5), .C(un14lto4), .Y(N_385));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[1]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[1]), .C(GND_net_1), .D(
        GND_net_1), .FCI(TC_Error_Counter_s_367_FCO), .S(
        \TC_Error_Counter_s[1] ), .Y(), .FCO(
        \TC_Error_Counter_cry[1]_net_1 ));
    CFG4 #( .INIT(16'h3F15) )  \Shift_reg_RNO_0[51]  (.A(N_349_1), .B(
        un1_TC_Packet_Counter17_5_net_1), .C(\State1[0]_net_1 ), .D(
        N_1463_mux), .Y(N_4558_i_1));
    CFG4 #( .INIT(16'h0800) )  Shift_reg_68_26_1580_i_i_N_6L11_RNO (.A(
        Shift_m3_2_1), .B(N_94_i), .C(Shift_reg_68_sn_N_56), .D(
        Shift_reg_1_sqmuxa_1_i_o3_0_o2_RNIJK1N_0_net_1), .Y(
        Shift_m3_2_3));
    SLE \TC_Packet_Counter[10]  (.D(\TC_Packet_Counter_s[10] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[10]));
    CFG3 #( .INIT(8'h57) )  \State1_ns_0_o2_0[0]  (.A(
        \block_counter[2]_net_1 ), .B(\block_counter[1]_net_1 ), .C(
        \block_counter[0]_net_1 ), .Y(TC_Packet_Counter17_i_0));
    CFG4 #( .INIT(16'hF0FB) )  Shift_reg_68_63_697_i_i_N_5L8 (.A(
        Shift_reg_68_1_2300_i_0_o2), .B(Shift_m4_e_1_sx), .C(
        Shift_reg_68_63_697_i_i_N_5L8_sx_net_1), .D(Shift_m8_i_a3_0_sx)
        , .Y(Shift_reg_68_63_697_i_i_N_5L8_net_1));
    CFG3 #( .INIT(8'h6A) )  Shift_reg_68_36_1321_i_m4_RNO (.A(
        \Shift_reg[20]_net_1 ), .B(\un1_Syn_reg[6] ), .C(N_1435), .Y(
        N_1433_mux));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_9_314_a2 (.A(CCA_NIRQ_c), .B(
        \Start_Buff[6]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3062));
    CFG4 #( .INIT(16'hFFFB) )  Shift_reg_68_24_1637_i_0_o2 (.A(N_55), 
        .B(un14lto4), .C(N_57), .D(N_265), .Y(N_62));
    CFG4 #( .INIT(16'h0880) )  Shift_reg_68_24_1637_i_0_a3_1_0 (.A(
        Shift_reg_68_50_5), .B(Shift_reg_68_sn_N_56), .C(
        \Shift_reg[39]_net_1 ), .D(N_398), .Y(
        Shift_reg_68_24_1637_i_0_a3_1_0_net_1));
    CFG3 #( .INIT(8'hD8) )  Shift_reg_68_4_2216_i_m4_bm (.A(
        Shift_reg_68_28_2_net_1), .B(RX_GPIO0_c), .C(
        \Shift_reg[47]_net_1 ), .Y(Shift_reg_68_4_2216_i_m4_bm_net_1));
    CFG4 #( .INIT(16'h78F0) )  Shift_reg_68_52_983_i_m4_am (.A(
        \Shift_reg_68_54_e_0[1] ), .B(Shift_reg_68_54_2), .C(
        \Shift_reg[2]_net_1 ), .D(\un1_Syn_reg[2] ), .Y(
        Shift_reg_68_52_983_i_m4_am_net_1));
    CFG2 #( .INIT(4'h4) )  un1_Syn_reg_67_1_x2_2_i_o3_RNIDKJK (.A(
        \un1_Syn_reg[0] ), .B(\State1[0]_net_1 ), .Y(
        Shift_reg_68_sn_N_16));
    SLE \TC_Error_Counter[9]  (.D(\TC_Error_Counter_s[9] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[9]));
    CFG4 #( .INIT(16'h0040) )  
        Shift_reg_68_0_2328_i_a7_0_0_a3_0_a3_0_a2_1_1_sx (.A(
        \un1_Syn_reg[0] ), .B(r_m1_e_1), .C(\un1_Syn_reg[4] ), .D(
        N_53_i), .Y(
        Shift_reg_68_0_2328_i_a7_0_0_a3_0_a3_0_a2_1_1_sx_net_1));
    CFG3 #( .INIT(8'h1B) )  Shift_reg_68_24_1637_i_0_0_N_2L1 (.A(N_62), 
        .B(RX_GPIO0_c), .C(\Shift_reg[39]_net_1 ), .Y(
        Shift_reg_68_24_1637_i_0_0_N_2L1_net_1));
    SLE \Shift_reg[41]  (.D(N_65), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[41]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  Shift_reg_68_30_1493_i_i (.A(N_114), .B(
        \Shift_reg[14]_net_1 ), .C(Shift_N_7_mux_0), .D(
        Shift_reg_68_30_1493_i_i_0_net_1), .Y(N_67));
    CFG3 #( .INIT(8'hFE) )  un1_block_counter (.A(
        \block_counter[2]_net_1 ), .B(\block_counter[1]_net_1 ), .C(
        \block_counter[0]_net_1 ), .Y(un1_block_counter_net_1));
    SLE \block_counter[0]  (.D(\block_counter_8[0]_net_1 ), .CLK(
        RX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \block_counter[0]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_34_1379_i_m4_ns (.A(
        Shift_reg_68_34_1379_i_m4_am_net_1), .B(
        Shift_reg_68_34_1379_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3960));
    CFG3 #( .INIT(8'hBA) )  Shift_reg_68_57_866_i_i_0_RNO (.A(
        Shift_m8_i_a3_0_sx_0), .B(Shift_reg_68_1_2300_i_0_o2), .C(
        Shift_m4_e_1_sx), .Y(Shift_m8_i_a3_0));
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_3_2244_i_m4_bm (.A(
        Shift_reg_68_28_1_1_net_1), .B(N_86), .C(RX_GPIO0_c), .D(
        \Shift_reg[46]_net_1 ), .Y(Shift_reg_68_3_2244_i_m4_bm_net_1));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_28_24_0_a3 (.A(
        \Bit_Counter[1]_net_1 ), .B(un14lto4), .C(un14lto5), .Y(
        Shift_reg_68_28_25_4));
    CFG4 #( .INIT(16'h1230) )  \block_counter_8[2]  (.A(CO0), .B(
        \un1_block_counter_7[0] ), .C(\block_counter[2]_net_1 ), .D(
        \block_counter[1]_net_1 ), .Y(\block_counter_8[2]_net_1 ));
    CFG3 #( .INIT(8'h6A) )  Shift_reg_68_27_1552_i_m4_am (.A(
        \Shift_reg[42]_net_1 ), .B(\un1_Syn_reg[5] ), .C(N_1461), .Y(
        Shift_reg_68_27_1552_i_m4_am_net_1));
    CFG4 #( .INIT(16'h0AFC) )  DataO_10_iv_0_0_RNO_24 (.A(
        \Shift_reg[55]_net_1 ), .B(\Shift_reg[51]_net_1 ), .C(
        \Shift_Bit_Counter[5]_net_1 ), .D(DataO_6_3_i_m2_1_2), .Y(
        N_339));
    CFG4 #( .INIT(16'h88B8) )  un1_Syn_reg_2_0_a3_1_RNI8JF3 (.A(
        \un1_Syn_reg[5] ), .B(\un1_Syn_reg[6] ), .C(N_244_2), .D(
        \un1_Syn_reg[2] ), .Y(Shift_reg_68_sn_m37_u_i_0));
    CFG4 #( .INIT(16'h2637) )  DataO_10_iv_0_0_RNO_1 (.A(
        \Shift_Bit_Counter[3]_net_1 ), .B(\Shift_Bit_Counter[4]_net_1 )
        , .C(N_2659), .D(N_2644), .Y(DataO_6_55_i_m2_1_2));
    CFG3 #( .INIT(8'hD8) )  \Shift_reg_68_28[34]  (.A(
        Shift_reg_68_28_16_net_1), .B(RX_GPIO0_c), .C(
        \Shift_reg[34]_net_1 ), .Y(N_104));
    CFG4 #( .INIT(16'hCC9C) )  \Shift_reg_RNO_0[13]  (.A(
        \un1_Syn_reg[2] ), .B(\Shift_reg[13]_net_1 ), .C(
        Shift_reg_68_50_2), .D(N_298), .Y(N_1451_mux));
    CFG4 #( .INIT(16'hB931) )  DataO_10_iv_0_0_RNO_11 (.A(
        \un22_DataO_i[2] ), .B(DataO_6_25_i_m3_1_2), .C(
        \Shift_reg[2]_net_1 ), .D(\Shift_reg[34]_net_1 ), .Y(N_400));
    CFG4 #( .INIT(16'h0015) )  \Shift_reg_RNO_1[13]  (.A(N_4080), .B(
        un1_TC_Packet_Counter17_5_net_1), .C(\State1[0]_net_1 ), .D(
        Shift_reg_68_29_1522_i_0_net_1), .Y(N_4079_i_1));
    CFG4 #( .INIT(16'h0800) )  Shift_reg_68_28_16_0 (.A(
        \Bit_Counter[2]_net_1 ), .B(un14lto4), .C(N_57), .D(un14lto0), 
        .Y(Shift_reg_68_28_42_4));
    SLE \Shift_reg[29]  (.D(N_4414_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[29]_net_1 ));
    CFG4 #( .INIT(16'hA008) )  Shift_reg_68_sn_m59_i_x3_RNI3Q7P3 (.A(
        N_54_i), .B(N_404), .C(\un1_Syn_reg[0] ), .D(
        Shift_reg_68_sn_N_9), .Y(
        Shift_reg_68_sn_m59_i_x3_RNI3Q7P3_net_1));
    CFG3 #( .INIT(8'h47) )  Shift_reg_68_63_697_i_i_N_5L8_sx (.A(
        Shift_reg_68_63_697_i_i_a2_0), .B(N_82), .C(
        Shift_reg_68_63_697_i_i_a2_0_0_net_1), .Y(
        Shift_reg_68_63_697_i_i_N_5L8_sx_net_1));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_3_2244_i_m4_ns (.A(
        Shift_reg_68_3_2244_i_m4_am_net_1), .B(
        Shift_reg_68_3_2244_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4680));
    CFG4 #( .INIT(16'h7FFF) )  un1_DataI_0_a3_a_a_a_a_a_a_sx (.A(
        un1_DataI_0_a3_a_a_a_a_a_a_N_3L3_net_1), .B(
        un1_DataI_0_a3_a_a_a_a_a_a_0_32), .C(
        un1_DataI_0_a3_a_a_a_a_a_a_N_2L1_net_1), .D(
        un1_DataI_0_a3_a_a_a_a_a_a_0_34), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_sx_net_1));
    CFG4 #( .INIT(16'h6996) )  Shift_reg_68_sn_m59_i_x3 (.A(
        \Syn_reg[4]_net_1 ), .B(\Parity[4]_net_1 ), .C(
        \Syn_reg[5]_net_1 ), .D(\Parity[5]_net_1 ), .Y(N_54_i));
    SLE \Start_Buff[6]  (.D(N_3072), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[6]_net_1 ));
    CFG4 #( .INIT(16'h0400) )  Shift_reg_68_38_1263_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_92_0)
        , .D(N_82), .Y(N_3868));
    CFG2 #( .INIT(4'hE) )  Shift_reg_68_28_21_a2_0_o2 (.A(un14lto0), 
        .B(\Bit_Counter[1]_net_1 ), .Y(N_265));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_10_2040_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_82), 
        .D(N_123_0), .Y(N_4516));
    SLE \TC_Packet_Counter[28]  (.D(\TC_Packet_Counter_s[28] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[28]));
    CFG2 #( .INIT(4'h4) )  \Syn_reg_RNO[3]  (.A(N_54), .B(
        \Syn_reg[2]_net_1 ), .Y(N_3287_i_0));
    SLE \Start_Sequence_counter[1]  (.D(
        \Start_Sequence_counter_9[1]_net_1 ), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\un6_DataO_i[1] ));
    CFG4 #( .INIT(16'h0080) )  \Parity_RNO[2]  (.A(CCA_NIRQ_c), .B(
        TC_Packet_Counter17_i_0), .C(N_3190), .D(N_277), .Y(N_3187_i_0)
        );
    SLE \Shift_reg[22]  (.D(N_3863_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[22]_net_1 ));
    CFG4 #( .INIT(16'hFCF5) )  Shift_reg_68_11_2010_i_2 (.A(
        \Shift_reg[54]_net_1 ), .B(Shift_reg_68_11_2010_i_a7_1_0_net_1)
        , .C(Shift_reg_68_11_2010_i_0_net_1), .D(
        Shift_reg_68_sn_N_84_mux), .Y(Shift_reg_68_11_2010_i_2_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIQEJ41[0]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[0]), .C(GND_net_1), .D(
        GND_net_1), .FCI(TC_Packet_Counter_cry_cy), .S(
        \TC_Packet_Counter_s[0] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[0] ));
    SLE \TC_Packet_Counter[14]  (.D(\TC_Packet_Counter_s[14] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[14]));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNILI5E6[17]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[17]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[16] ), .S(
        \TC_Packet_Counter_s[17] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[17] ));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[45]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4705), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4702_i_0));
    CFG3 #( .INIT(8'h20) )  Shift_reg_68_28_15_0 (.A(
        \Bit_Counter[2]_net_1 ), .B(N_374), .C(un14lto4), .Y(
        Shift_reg_68_28_41_4));
    CFG4 #( .INIT(16'hDF8A) )  \un1_block_counter_3[0]  (.A(CCA_NIRQ_c)
        , .B(\State2[0]_net_1 ), .C(\State2[1]_net_1 ), .D(
        un1_block_counter_net_1), .Y(Shift_Bit_Countere));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_s[31]  (.A(VCC_net_1)
        , .B(CLTU_0_TC_Error_Counter[31]), .C(GND_net_1), .D(GND_net_1)
        , .FCI(\TC_Error_Counter_cry[30]_net_1 ), .S(
        \TC_Error_Counter_s[31]_net_1 ), .Y(), .FCO());
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_12_1982_i_m4_bm (.A(
        Shift_reg_68_28_10_1_net_1), .B(N_57), .C(RX_GPIO0_c), .D(
        \Shift_reg[55]_net_1 ), .Y(Shift_reg_68_12_1982_i_m4_bm_net_1));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_sn_m23_0_a2_RNI3IHS (.A(
        Shift_reg_68_sn_N_24), .B(\un1_Syn_reg[0] ), .C(
        \un1_Syn_reg[6] ), .Y(\Shift_reg_68_54_e_0[1] ));
    CFG4 #( .INIT(16'h2367) )  DataO_10_iv_0_0_RNO_15 (.A(
        \un22_DataO_i[0] ), .B(\un22_DataO_i[1] ), .C(N_339), .D(N_333)
        , .Y(DataO_6_15_1_2));
    CFG4 #( .INIT(16'h3F15) )  \Shift_reg_RNO_0[5]  (.A(N_349_1), .B(
        un1_TC_Packet_Counter17_5_net_1), .C(\State1[0]_net_1 ), .D(
        N_1438_mux), .Y(N_3558_i_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIO5CV6[20]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[20]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[19] ), .S(
        \TC_Packet_Counter_s[20] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[20] ));
    CFG4 #( .INIT(16'h6996) )  Shift_reg_68_sn_m21_0_a2_0_x2 (.A(
        \Parity[1]_net_1 ), .B(\Syn_reg[1]_net_1 ), .C(
        \Syn_reg[6]_net_1 ), .D(\Parity[6]_net_1 ), .Y(N_97_i));
    CFG4 #( .INIT(16'hFFF8) )  Shift_reg_68_57_866_i_i (.A(N_114), .B(
        \Shift_reg[6]_net_1 ), .C(Shift_N_10_mux), .D(
        Shift_reg_68_57_866_i_i_0_net_1), .Y(N_71));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[7]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[7]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[6]_net_1 ), .S(
        \TC_Error_Counter_s[7] ), .Y(), .FCO(
        \TC_Error_Counter_cry[7]_net_1 ));
    SLE \TC_Packet_Counter[13]  (.D(\TC_Packet_Counter_s[13] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[13]));
    CFG4 #( .INIT(16'hCCCD) )  Shift_reg_68_1_2300_i_0_0 (.A(N_86), .B(
        N_74), .C(RX_GPIO0_c), .D(Shift_reg_68_1_2300_i_0_o3_1_0_net_1)
        , .Y(Shift_reg_68_1_2300_i_0_0_net_1));
    CFG2 #( .INIT(4'hB) )  Parity_16_2_480_i_0_o2_0 (.A(
        \Parity_Counter[1]_net_1 ), .B(\Parity_Counter[2]_net_1 ), .Y(
        Parity_16_3_456_i_o4_0));
    CFG4 #( .INIT(16'h0048) )  un1_Syn_reg_67_1_a6_3 (.A(
        \un1_Syn_reg[6] ), .B(un1_Syn_reg_67_1_a6_3_0_net_1), .C(
        \un1_Syn_reg[5] ), .D(N_53_i), .Y(N_2847));
    CFG2 #( .INIT(4'h1) )  Shift_reg_68_28_51_0 (.A(N_265), .B(N_34), 
        .Y(Shift_reg_68_28_51_0_net_1));
    CFG3 #( .INIT(8'h02) )  Shift_reg_68_28_22_1 (.A(
        \Bit_Counter[3]_net_1 ), .B(un14lto4), .C(un14lto5), .Y(
        Shift_reg_68_28_22_1_net_1));
    SLE \TC_Packet_Counter[3]  (.D(\TC_Packet_Counter_s[3] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[3]));
    CFG3 #( .INIT(8'h41) )  \Start_Sequence_counter_9[0]  (.A(
        \un1_block_counter_7[0] ), .B(\un6_DataO_i[0] ), .C(
        un1_DataO41_18), .Y(\Start_Sequence_counter_9[0]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \Syn_reg_RNO[1]  (.A(N_54), .B(
        \Syn_reg[0]_net_1 ), .Y(N_3319_i_0));
    SLE \Start_Buff[12]  (.D(Start_Buff_10_14_259_a2_net_1), .CLK(
        RX_GPIO1_c), .EN(un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[12]_net_1 ));
    CFG4 #( .INIT(16'h23EF) )  Shift_reg_68_19_1783_i_0_o3 (.A(N_381), 
        .B(Shift_reg_68_sn_N_84_mux), .C(\un1_Syn_reg[0] ), .D(N_287), 
        .Y(N_388));
    CFG4 #( .INIT(16'h78F0) )  \Shift_reg_RNO_1[5]  (.A(
        \un1_Syn_reg[0] ), .B(Shift_reg_68_50_net_1), .C(
        \Shift_reg[5]_net_1 ), .D(\un1_Syn_reg[5] ), .Y(N_1438_mux));
    CFG4 #( .INIT(16'h3337) )  Shift_reg_68_38_1263_i_0 (.A(
        \Shift_reg[22]_net_1 ), .B(CCA_NIRQ_c), .C(
        Shift_reg_68_sn_N_56), .D(N_82), .Y(N_3863_i_1_1));
    SLE \TC_Packet_Counter[0]  (.D(\TC_Packet_Counter_s[0] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[0]));
    CFG3 #( .INIT(8'h10) )  \Shift_reg_RNO[51]  (.A(N_346), .B(
        Shift_reg_68_8_2099_i_0_1_net_1), .C(N_4558_i_1), .Y(
        N_4558_i_0));
    SLE \Shift_reg[30]  (.D(N_4389_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[30]_net_1 ));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[40]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4154), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4151_i_0));
    CFG4 #( .INIT(16'hFBFF) )  Shift_reg_68_30_1493_i_i_o3_1 (.A(
        \Bit_Counter[2]_net_1 ), .B(\Bit_Counter[3]_net_1 ), .C(N_57), 
        .D(un14lto0), .Y(N_210));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNISPDD8[28]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[28]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[27] ), .S(
        \TC_Packet_Counter_s[28] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[28] ));
    CFG3 #( .INIT(8'h10) )  Shift_reg_68_28_28_1 (.A(
        \Bit_Counter[3]_net_1 ), .B(un14lto4), .C(un14lto5), .Y(
        Shift_reg_68_28_28_1_net_1));
    CFG4 #( .INIT(16'h6C80) )  Shift_reg_68_50_1 (.A(\un1_Syn_reg[2] ), 
        .B(N_53_i), .C(\un1_Syn_reg[0] ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_50_5));
    CFG4 #( .INIT(16'hF078) )  Shift_reg_68_34_1379_i_m4_am (.A(
        \Shift_reg_68_54_e_0[4] ), .B(Shift_reg_68_54_net_1), .C(
        \Shift_reg[18]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_34_1379_i_m4_am_net_1));
    CFG4 #( .INIT(16'hA202) )  Shift_reg_68_26_1580_i_i_1_tz (.A(
        \Shift_reg[41]_net_1 ), .B(N_53_i), .C(N_82), .D(N_219), .Y(
        Shift_reg_68_26_1580_i_i_1_tz_net_1));
    SLE \Shift_reg[19]  (.D(N_3935_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[19]_net_1 ));
    SLE \Shift_reg[2]  (.D(N_3627_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[2]_net_1 ));
    SLE \TC_Packet_Counter[30]  (.D(\TC_Packet_Counter_s[30] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[30]));
    CFG4 #( .INIT(16'h0080) )  Shift_reg_68_37_1293_i_0_a2_2_1 (.A(
        \Shift_reg[21]_net_1 ), .B(\un1_Syn_reg[0] ), .C(
        \un1_Syn_reg[6] ), .D(N_381), .Y(
        Shift_reg_68_37_1293_i_0_a2_2_1_net_1));
    SLE \block_counter[2]  (.D(\block_counter_8[2]_net_1 ), .CLK(
        RX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \block_counter[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  Start_Buff_10_2_391_a2_1 (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .Y(N_2992));
    SLE \Syn_reg[3]  (.D(N_3287_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_15_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Syn_reg[3]_net_1 ));
    CFG2 #( .INIT(4'h2) )  Shift_reg_68_57_866_i_i_a2_3_1_1 (.A(
        Shift_reg_1_sqmuxa_1_i_o3_0_o2_RNIJK1N_0_net_1), .B(
        Shift_reg_68_1_2300_i_0_o2), .Y(
        Shift_reg_68_57_866_i_i_a2_3_1_1_net_1));
    CFG4 #( .INIT(16'h0020) )  un1_Start_Buff_1_5 (.A(
        \Start_Buff[13]_net_1 ), .B(\Start_Buff[12]_net_1 ), .C(
        \Start_Buff[11]_net_1 ), .D(\Start_Buff[10]_net_1 ), .Y(
        un1_Start_Buff_1_5_0));
    CFG4 #( .INIT(16'h0084) )  un1_Syn_reg_67_1_a6_2 (.A(
        \un1_Syn_reg[6] ), .B(un1_Syn_reg_67_1_a6_2_1_net_1), .C(
        \un1_Syn_reg[5] ), .D(N_53_i), .Y(N_2846));
    SLE \TC_Packet_Counter[6]  (.D(\TC_Packet_Counter_s[6] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[6]));
    SLE \Shift_reg[12]  (.D(N_75), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[12]_net_1 ));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_679_a2 (.A(CCA_NIRQ_c), .B(
        \Start_Buff[12]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3366));
    SLE \Shift_reg[26]  (.D(N_3767_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[26]_net_1 ));
    CFG3 #( .INIT(8'h80) )  un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_x_RNO (.A(
        \Shift_reg[42]_net_1 ), .B(\Shift_reg[48]_net_1 ), .C(
        \Shift_reg[47]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_x_RNO_net_1));
    CFG4 #( .INIT(16'h0020) )  Shift_reg_68_13_1953_i_i_N_4L5_N_5L8 (
        .A(Shift_reg_1_sqmuxa_1_i_o3_0_o2_RNIJK1N_0_net_1), .B(
        Shift_reg_68_sn_N_56), .C(
        Shift_reg_68_13_1953_i_i_N_4L5_N_3L4_net_1), .D(
        Shift_reg_68_1_2300_i_0_o2), .Y(
        Shift_reg_68_13_1953_i_i_N_4L5_N_5L8_net_1));
    SLE \Shift_reg[28]  (.D(N_61), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[28]_net_1 ));
    CFG4 #( .INIT(16'h2367) )  DataO_10_iv_0_0_RNO_19 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[38]_net_1 ), .D(\Shift_reg[6]_net_1 ), .Y(
        DataO_6_25_i_m3_1_2));
    CFG4 #( .INIT(16'hB3FF) )  Shift_reg_1_sqmuxa_1_i_o3_0 (.A(
        un14lto5), .B(\State1[0]_net_1 ), .C(N_436_1), .D(
        TC_Packet_Counter17_i_0), .Y(N_57));
    CFG4 #( .INIT(16'hFEEE) )  Shift_reg_68_21_1723_i_i_3 (.A(
        Shift_reg_68_21_1723_i_i_3_1), .B(N_227), .C(
        \Shift_reg[36]_net_1 ), .D(N_250), .Y(N_56));
    CFG4 #( .INIT(16'hFBFF) )  Shift_reg_68_46_1115_i_i_N_8L17 (.A(
        Shift_reg_68_1_2300_i_0_o2), .B(\Shift_reg[27]_net_1 ), .C(
        Shift_reg_68_46_1115_i_i_N_8L17_1_net_1), .D(N_215), .Y(
        Shift_reg_68_46_1115_i_i_N_8L17_net_1));
    CFG4 #( .INIT(16'h0080) )  un1_DataI_0_a3_a_a_a_a_a_a_N_3L3 (.A(
        RX_GPIO0_c), .B(\Shift_reg[39]_net_1 ), .C(
        \Shift_reg[34]_net_1 ), .D(\Shift_reg[12]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_N_3L3_net_1));
    SLE \TC_Packet_Counter[2]  (.D(\TC_Packet_Counter_s[2] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[2]));
    CFG4 #( .INIT(16'h0015) )  \Shift_reg_RNO_1[23]  (.A(N_3842), .B(
        un1_TC_Packet_Counter17_5_net_1), .C(\State1[0]_net_1 ), .D(
        Shift_reg_68_39_1233_i_0_net_1), .Y(N_3841_i_1));
    CFG3 #( .INIT(8'hCE) )  Shift_reg_1_sqmuxa_1_i_o3_0_o2_RNIJK1N (.A(
        \State1[0]_net_1 ), .B(\un1_Syn_reg[0] ), .C(N_58), .Y(N_82));
    CFG2 #( .INIT(4'h8) )  Block_ErrO_2_sqmuxa_1_i_a0_0 (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .Y(
        Block_ErrO_2_sqmuxa_1_i_a1_0));
    CFG3 #( .INIT(8'h02) )  Shift_reg_68_28_35_1 (.A(un14lto5), .B(
        N_265), .C(N_387), .Y(Shift_reg_68_28_35_1_net_1));
    CFG4 #( .INIT(16'h3705) )  Shift_reg_68_30_1493_i_i_0 (.A(N_74), 
        .B(Shift_N_5), .C(Shift_N_9_0), .D(Shift_m2_0_3), .Y(
        Shift_reg_68_30_1493_i_i_0_net_1));
    CFG4 #( .INIT(16'h3F15) )  \Shift_reg_RNO_0[15]  (.A(N_349_1), .B(
        un1_TC_Packet_Counter17_5_net_1), .C(\State1[0]_net_1 ), .D(
        N_1472_mux), .Y(N_4032_i_1));
    CFG2 #( .INIT(4'h8) )  Shift_reg_68_sn_m57_i_o3_RNISOJH (.A(
        \un1_Syn_reg[0] ), .B(\un1_Syn_reg[5] ), .Y(
        \Shift_reg_68_54_e_0[29] ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIINCM7[24]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[24]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[23] ), .S(
        \TC_Packet_Counter_s[24] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[24] ));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_12_281_a2 (.A(CCA_NIRQ_c), 
        .B(\Start_Buff[9]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3032));
    CFG4 #( .INIT(16'hF078) )  \Shift_reg_RNO_1[15]  (.A(
        \un1_Syn_reg[0] ), .B(Shift_reg_68_50_net_1), .C(
        \Shift_reg[15]_net_1 ), .D(\un1_Syn_reg[5] ), .Y(N_1472_mux));
    CFG3 #( .INIT(8'h40) )  Shift_reg_68_28_10_1 (.A(un14lto0), .B(
        Shift_reg_68_28_9_2), .C(Shift_reg_68_28_6_4), .Y(
        Shift_reg_68_28_10_1_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIEEKI4[8]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[8]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Packet_Counter_cry[7] ), .S(
        \TC_Packet_Counter_s[8] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[8] ));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[26]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3770), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3767_i_0));
    CFG4 #( .INIT(16'hFBC8) )  Shift_reg_68_9_2070_i_0_m2 (.A(N_86), 
        .B(N_82), .C(Shift_reg_68_9_2070_i_0_o2_1_1_net_1), .D(N_268), 
        .Y(N_81));
    SLE \Syn_reg[4]  (.D(N_3275_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_15_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Syn_reg[4]_net_1 ));
    CFG4 #( .INIT(16'h5D0C) )  Shift_reg_68_46_1115_i_i_N_9L19 (.A(
        Shift_reg_68_46_1115_i_i_N_8L17_net_1), .B(N_253), .C(N_215), 
        .D(Shift_reg_68_sn_N_84_mux), .Y(Shift_reg_68_46_1115_i_i_1));
    SLE \Shift_reg[49]  (.D(N_59), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[49]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  \State1_ns_0_a5_2_9[0]  (.A(
        \Start_Buff[12]_net_1 ), .B(\State1[0]_net_1 ), .C(
        \State1_ns_0_a5_2_4[0]_net_1 ), .D(\State1_ns_0_a5_2_6[0] ), 
        .Y(\State1_ns_0_a5_2_9[0]_net_1 ));
    CFG4 #( .INIT(16'hF99F) )  \Syn_reg_RNIUMFH1[3]  (.A(
        \Syn_reg[3]_net_1 ), .B(\Parity[3]_net_1 ), .C(
        \Syn_reg[2]_net_1 ), .D(\Parity[2]_net_1 ), .Y(N_404));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[17]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3985), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3982_i_0));
    CFG4 #( .INIT(16'h0060) )  Shift_reg_68_10_2040_i_a7_1_RNO (.A(
        \un1_Syn_reg[2] ), .B(N_53_i), .C(\un1_Syn_reg[0] ), .D(
        \un1_Syn_reg[6] ), .Y(N_1463));
    CFG3 #( .INIT(8'hE4) )  \un1_block_counter_7_ns[0]  (.A(CCA_NIRQ_c)
        , .B(\un1_block_counter_7_am[0]_net_1 ), .C(
        \un1_block_counter_7_bm[0]_net_1 ), .Y(
        \un1_block_counter_7[0] ));
    CFG4 #( .INIT(16'h2112) )  \Syn_reg_RNO[2]  (.A(\Syn_reg[6]_net_1 )
        , .B(N_54), .C(RX_GPIO0_c), .D(\Syn_reg[1]_net_1 ), .Y(
        N_3301_i_0));
    CFG4 #( .INIT(16'h0001) )  \Shift_reg_RNI1EJ6[33]  (.A(
        \Shift_reg[36]_net_1 ), .B(\Shift_reg[33]_net_1 ), .C(
        \Shift_reg[28]_net_1 ), .D(\Shift_reg[35]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_44));
    CFG3 #( .INIT(8'hD8) )  Shift_reg_68_58_838_i_m4_bm (.A(
        Shift_reg_68_28_47_net_1), .B(RX_GPIO0_c), .C(
        \Shift_reg[7]_net_1 ), .Y(Shift_reg_68_58_838_i_m4_bm_net_1));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_17_1839_i_a7_2 (.A(
        Shift_reg_68_sn_N_56), .B(\Shift_reg[32]_net_1 ), .C(N_82), .Y(
        N_4346));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[22]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[22]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[21]_net_1 ), .S(
        \TC_Error_Counter_s[22] ), .Y(), .FCO(
        \TC_Error_Counter_cry[22]_net_1 ));
    CFG4 #( .INIT(16'hF078) )  Shift_reg_68_59_810_i_m4_am (.A(
        \Shift_reg_68_54_e_0[8] ), .B(Shift_reg_68_54_2), .C(
        \Shift_reg[8]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_59_810_i_m4_am_net_1));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[4]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3583), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3580_i_0));
    SLE \TC_Error_Counter[24]  (.D(\TC_Error_Counter_s[24] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[24]));
    SLE \Shift_Bit_Counter[5]  (.D(\Shift_Bit_Counter_s[5]_net_1 ), 
        .CLK(RX_GPIO1_c), .EN(Shift_Bit_Countere), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_Bit_Counter[5]_net_1 ));
    SLE \Shift_reg[42]  (.D(N_4101_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[42]_net_1 ));
    CFG4 #( .INIT(16'h8068) )  Shift_reg_68_50_0 (.A(\un1_Syn_reg[2] ), 
        .B(N_53_i), .C(\un1_Syn_reg[0] ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_50_9));
    CFG3 #( .INIT(8'hDF) )  \Shift_reg_68_38_i_o3[39]  (.A(
        \un1_Syn_reg[6] ), .B(N_53_i), .C(\un1_Syn_reg[0] ), .Y(N_398));
    CFG4 #( .INIT(16'h0AFC) )  DataO_10_iv_0_0_RNO_4 (.A(
        \Shift_reg[44]_net_1 ), .B(\Shift_reg[40]_net_1 ), .C(
        \Shift_Bit_Counter[5]_net_1 ), .D(DataO_6_44_1_2), .Y(N_2673));
    CFG2 #( .INIT(4'h2) )  Shift_reg_68_28_6_0 (.A(Shift_reg_68_28_6_4)
        , .B(N_265), .Y(Shift_reg_68_28_6_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[14]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[14]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[13]_net_1 ), .S(
        \TC_Error_Counter_s[14] ), .Y(), .FCO(
        \TC_Error_Counter_cry[14]_net_1 ));
    CFG4 #( .INIT(16'h78F0) )  Shift_reg_68_40_1205_i_m4_am (.A(
        Shift_reg_68_43_2), .B(Shift_reg_68_54_4), .C(
        \Shift_reg[24]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_40_1205_i_m4_am_net_1));
    CFG4 #( .INIT(16'h4000) )  Shift_reg_68_28_29_1 (.A(un14lto4), .B(
        \Bit_Counter[2]_net_1 ), .C(un14lto5), .D(Shift_reg_68_28_29_3)
        , .Y(Shift_reg_68_28_29_1_net_1));
    CFG4 #( .INIT(16'h0080) )  \Shift_reg_RNO[43]  (.A(N_4752_i_1), .B(
        \Shift_reg_RNO_1[43]_net_1 ), .C(CCA_NIRQ_c), .D(N_4756), .Y(
        N_4752_i_0));
    CFG4 #( .INIT(16'h80A0) )  Shift_reg_68_35_1349_i_a7_1_1 (.A(
        \State1[0]_net_1 ), .B(un1_TC_Packet_Counter17_3_net_1), .C(
        Shift_reg_68_sn_N_56), .D(Shift_reg_68_sn_N_73), .Y(N_349_1));
    CFG4 #( .INIT(16'h000D) )  un1_DataO41_22_0_a3_0_4_RNIRAVS (.A(
        un1_DataO41_22_0_a3_0_3_net_1), .B(
        un1_TC_Packet_Counter17_3_net_1), .C(un1_DataO41_22_0_0_net_1), 
        .D(un1_DataO41_22_0_1_net_1), .Y(un1_DataO41_22_i_0));
    CFG3 #( .INIT(8'h08) )  Shift_reg_68_28_25_0 (.A(
        Shift_reg_68_28_25_4), .B(\Bit_Counter[3]_net_1 ), .C(un14lto0)
        , .Y(Shift_reg_68_28_25_0_net_1));
    CFG3 #( .INIT(8'hAC) )  Shift_reg_68_sn_m59_i_x3_RNI4Q8U2 (.A(
        Shift_reg_68_sn_m59_i_x3_RNI590H_net_1), .B(
        Shift_reg_68_sn_m72_6_am_1), .C(N_1431), .Y(N_2548));
    CFG3 #( .INIT(8'h10) )  \Parity_RNO[3]  (.A(N_2969_1), .B(N_277), 
        .C(N_78), .Y(N_3167_i_0));
    CFG4 #( .INIT(16'h0060) )  un1_Syn_reg_67_1_a6_3_0 (.A(
        \Parity[0]_net_1 ), .B(\Syn_reg[0]_net_1 ), .C(N_376), .D(
        \un1_Syn_reg[4] ), .Y(un1_Syn_reg_67_1_a6_3_0_net_1));
    CFG4 #( .INIT(16'hFE10) )  Parity_16_1_505_i_0_m2 (.A(
        \Parity_Counter[0]_net_1 ), .B(Parity_16_1_505_i_0_o2_0_net_1), 
        .C(RX_GPIO0_c), .D(\Parity[0]_net_1 ), .Y(N_275));
    CFG2 #( .INIT(4'h2) )  Shift_reg_68_sn_m57_i_o3_RNISOJH_1 (.A(
        \un1_Syn_reg[0] ), .B(\un1_Syn_reg[5] ), .Y(
        \Shift_reg_68_54_e_0[10] ));
    SLE \Shift_reg[16]  (.D(N_4007_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[16]_net_1 ));
    CFG3 #( .INIT(8'h10) )  Shift_reg_68_30_1493_i_i_RNO (.A(N_102), 
        .B(N_210), .C(N_253), .Y(Shift_N_7_mux_0));
    CFG4 #( .INIT(16'h4567) )  DataO_10_iv_0_0_RNO_12 (.A(
        \un22_DataO_i[1] ), .B(\un22_DataO_i[0] ), .C(N_325), .D(N_322)
        , .Y(DataO_6_30_1_2));
    SLE \TC_Error_Counter[13]  (.D(\TC_Error_Counter_s[13] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[13]));
    SLE \Shift_reg[18]  (.D(N_3957_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[18]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \Bit_Counter_cry[4]  (.A(VCC_net_1), 
        .B(un14lto4), .C(GND_net_1), .D(GND_net_1), .FCI(
        \Bit_Counter_cry[3]_net_1 ), .S(\Bit_Counter_s[4] ), .Y(), 
        .FCO(\Bit_Counter_cry[4]_net_1 ));
    CFG3 #( .INIT(8'h20) )  Shift_reg_1_sqmuxa_1_i_o3_0_o2_RNIJK1N_0 (
        .A(\State1[0]_net_1 ), .B(\un1_Syn_reg[0] ), .C(N_58), .Y(
        Shift_reg_1_sqmuxa_1_i_o3_0_o2_RNIJK1N_0_net_1));
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_34_1379_i_m4_bm (.A(
        Shift_reg_68_28_30_0_net_1), .B(N_86), .C(RX_GPIO0_c), .D(
        \Shift_reg[18]_net_1 ), .Y(Shift_reg_68_34_1379_i_m4_bm_net_1));
    CFG4 #( .INIT(16'h78F0) )  Shift_reg_68_14_1925_i_m4_am (.A(
        \Shift_reg_68_54_e_0[29] ), .B(Shift_reg_68_54_4), .C(
        \Shift_reg[29]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_14_1925_i_m4_am_net_1));
    CFG3 #( .INIT(8'h04) )  Shift_reg_68_63_697_i_i_a2_2_1 (.A(N_87), 
        .B(N_253), .C(N_103), .Y(N_199_1));
    SLE \Shift_reg[9]  (.D(N_73), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[9]_net_1 ));
    CFG4 #( .INIT(16'h0080) )  un1_DataI_0_a3_a_a_a_a_a_a_x (.A(
        un1_DataI_0_a3_a_a_a_a_a_a_0_56), .B(
        un1_DataI_0_a3_a_a_a_a_a_a_0_58), .C(
        un1_DataI_0_a3_a_a_a_a_a_a_0_33), .D(
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_x_net_1), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_x_net_1));
    CFG4 #( .INIT(16'h7FFF) )  un1_DataI_0_a3_a_a_a_a_a_a_N_5L7 (.A(
        un1_DataI_0_a3_a_a_a_a_a_a_N_3L3_net_1), .B(
        un1_DataI_0_a3_a_a_a_a_a_a_0_32), .C(
        un1_DataI_0_a3_a_a_a_a_a_a_N_2L1_net_1), .D(
        un1_DataI_0_a3_a_a_a_a_a_a_0_34), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_N_5L7_net_1));
    CFG4 #( .INIT(16'hFFF9) )  Shift_reg_68_30_1493_i_i_o3_0 (.A(
        \Parity[6]_net_1 ), .B(\Syn_reg[6]_net_1 ), .C(
        \un1_Syn_reg[5] ), .D(N_53_i), .Y(N_122));
    CFG3 #( .INIT(8'h63) )  Shift_reg_68_12_1982_i_m4_am (.A(
        Shift_reg_68_sn_N_49), .B(N_1456_mux), .C(
        \Shift_reg_68_54_e_1[55] ), .Y(
        Shift_reg_68_12_1982_i_m4_am_net_1));
    CFG4 #( .INIT(16'h0007) )  \Shift_reg_RNO[35]  (.A(
        \State1[0]_net_1 ), .B(un1_TC_Packet_Counter17_5_net_1), .C(
        N_4275), .D(Shift_reg_68_20_1753_i_2_net_1), .Y(N_4270_i_0));
    CFG4 #( .INIT(16'h660A) )  \un1_Syn_reg_i_o3_RNI1C5B1[2]  (.A(
        N_53_i), .B(\un1_Syn_reg[2] ), .C(Shift_reg_68_sn_N_50), .D(
        \un1_Syn_reg[6] ), .Y(N_2188));
    CFG4 #( .INIT(16'h51EA) )  Shift_reg_68_12_1982_i_m4_am_RNO (.A(
        \State1[0]_net_1 ), .B(un1_Start_Buff_1_net_1), .C(RX_GPIO0_c), 
        .D(\Shift_reg[55]_net_1 ), .Y(N_1456_mux));
    CFG2 #( .INIT(4'hD) )  Parity_16_5_407_i_o4_0 (.A(
        \Parity_Counter[1]_net_1 ), .B(\Parity_Counter[2]_net_1 ), .Y(
        Parity_16_5_407_i_o4_0_net_1));
    CFG4 #( .INIT(16'hB931) )  DataO_10_iv_0_0_RNO_2 (.A(
        \un22_DataO_i[2] ), .B(DataO_6_41_i_m2_1_2), .C(
        \Shift_reg[10]_net_1 ), .D(\Shift_reg[42]_net_1 ), .Y(N_314));
    CFG4 #( .INIT(16'h0AFC) )  DataO_10_iv_0_0_RNO_21 (.A(
        \Shift_reg[37]_net_1 ), .B(\Shift_reg[33]_net_1 ), .C(
        \Shift_Bit_Counter[5]_net_1 ), .D(DataO_6_21_i_m2_1_2), .Y(
        N_322));
    CFG3 #( .INIT(8'h10) )  Shift_reg_68_28_11_0 (.A(
        \Bit_Counter[2]_net_1 ), .B(un14lto0), .C(N_436_1), .Y(
        Shift_reg_68_28_11_0_net_1));
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_33_1407_i_m4_bm (.A(
        Shift_reg_68_28_29_1_net_1), .B(N_374), .C(RX_GPIO0_c), .D(
        \Shift_reg[17]_net_1 ), .Y(Shift_reg_68_33_1407_i_m4_bm_net_1));
    CFG3 #( .INIT(8'hF7) )  Shift_reg_68_28_17_1_i_o2 (.A(
        \Bit_Counter[2]_net_1 ), .B(\State1[0]_net_1 ), .C(N_58), .Y(
        N_92));
    SLE \TC_Error_Counter[1]  (.D(\TC_Error_Counter_s[1] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[1]));
    CFG4 #( .INIT(16'h0020) )  un1_DataI_0_a3_a_a_a_a_a_a (.A(
        un1_DataI_0_a3_a_a_a_a_a_a_0_56), .B(
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_net_1), .C(
        un1_DataI_0_a3_a_a_a_a_a_a_0_58), .D(
        un1_DataI_0_a3_a_a_a_a_a_a_sx_net_1), .Y(un1_DataI));
    CFG3 #( .INIT(8'h10) )  Shift_reg_68_26_1580_i_i_N_4L6 (.A(N_57), 
        .B(N_91), .C(Shift_reg_68_26_1580_i_i_N_2L1_net_1), .Y(
        Shift_reg_68_26_1580_i_i_N_4L6_net_1));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_11_292_a2 (.A(CCA_NIRQ_c), 
        .B(\Start_Buff[8]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3042));
    CFG4 #( .INIT(16'h02A2) )  Shift_reg_1_sqmuxa_1_i_o3_0_RNIK3RB2 (
        .A(N_57), .B(N_2188), .C(\un1_Syn_reg[0] ), .D(
        Shift_reg_68_sn_N_82_mux), .Y(Shift_reg_68_sn_N_56));
    ARI1 #( .INIT(20'h48800) )  \Shift_Bit_Counter_cry[0]  (.A(
        VCC_net_1), .B(\un22_DataO_i[0] ), .C(
        \Shift_Bit_Counter_cry_cy_Y[0] ), .D(GND_net_1), .FCI(
        Shift_Bit_Counter_cry_cy), .S(\Shift_Bit_Counter_s[0] ), .Y(), 
        .FCO(\Shift_Bit_Counter_cry[0]_net_1 ));
    SLE \Shift_reg[6]  (.D(N_71), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[6]_net_1 ));
    CFG4 #( .INIT(16'hA600) )  Shift_reg_68_23_1667_i_i_a2_0 (.A(
        \Shift_reg[38]_net_1 ), .B(N_53_i), .C(N_101), .D(N_250), .Y(
        N_172));
    SLE \Parity[2]  (.D(N_3187_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_10_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Parity[2]_net_1 ));
    CFG2 #( .INIT(4'h7) )  Parity_16_4_431_i_0_o3 (.A(
        TC_Packet_Counter17_i_0), .B(CCA_NIRQ_c), .Y(N_2969_1));
    SLE \TC_Packet_Counter[12]  (.D(\TC_Packet_Counter_s[12] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[12]));
    CFG3 #( .INIT(8'h6F) )  Shift_reg_68_57_866_i_i_o3 (.A(
        \Parity[6]_net_1 ), .B(\Syn_reg[6]_net_1 ), .C(
        \un1_Syn_reg[2] ), .Y(N_123));
    CFG2 #( .INIT(4'h7) )  un1_State1_0 (.A(TC_Packet_Counter18_i_0), 
        .B(\State1[0]_net_1 ), .Y(un1_State1_0_net_1));
    CFG2 #( .INIT(4'h4) )  un1_DataO41_27_a1_0 (.A(N_277), .B(
        TC_Packet_Counter17_i_0), .Y(un1_DataO41_27_a1_0_net_1));
    CFG4 #( .INIT(16'h0010) )  Shift_reg_68_46_1115_i_i_N_8L17_1 (.A(
        un1_TC_Packet_Counter17_1_net_1), .B(un1_DataI), .C(
        Shift_m3_e_3), .D(\State1_ns_0_o5_2[0]_net_1 ), .Y(
        Shift_reg_68_46_1115_i_i_N_8L17_1_net_1));
    CFG2 #( .INIT(4'h4) )  Shift_reg_68_54_RNO (.A(
        Shift_reg_68_sn_N_32), .B(\State1[0]_net_1 ), .Y(
        Shift_reg_68_sn_N_33));
    CFG4 #( .INIT(16'h006C) )  \Start_Sequence_counter_9[2]  (.A(
        \un6_DataO_i[1] ), .B(\un6_DataO_i[2] ), .C(CO0_1), .D(
        \un1_block_counter_7[0] ), .Y(
        \Start_Sequence_counter_9[2]_net_1 ));
    CFG3 #( .INIT(8'h10) )  Shift_reg_68_28_45_0 (.A(
        \Bit_Counter[2]_net_1 ), .B(un14lto0), .C(N_21_i), .Y(
        Shift_reg_68_28_45_0_net_1));
    CFG4 #( .INIT(16'h5557) )  un1_TC_Packet_Counter17_5 (.A(
        TC_Packet_Counter17_i_0), .B(\State1_ns_0_o5_2[0]_net_1 ), .C(
        un1_TC_Packet_Counter17_3_net_1), .D(
        \State1_ns_0_o5_3[0]_net_1 ), .Y(
        un1_TC_Packet_Counter17_5_net_1));
    CFG4 #( .INIT(16'h0FAC) )  DataO_10_iv_0_0_RNO_25 (.A(
        \Shift_reg[53]_net_1 ), .B(\Shift_reg[49]_net_1 ), .C(
        DataO_6_6_i_m2_1_2), .D(\Shift_Bit_Counter[5]_net_1 ), .Y(
        N_333));
    CFG3 #( .INIT(8'hB3) )  Shift_reg_68_24_1637_i_0_a2_0 (.A(
        Shift_reg_68_sn_N_82_mux), .B(N_57), .C(\un1_Syn_reg[0] ), .Y(
        N_287));
    SLE \Shift_reg[46]  (.D(N_4677_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[46]_net_1 ));
    CFG3 #( .INIT(8'h6C) )  \Shift_reg_RNO_1[32]  (.A(
        Shift_reg_68_50_2), .B(\Shift_reg[32]_net_1 ), .C(N_53_i), .Y(
        N_1452_mux));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[30]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4392), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4389_i_0));
    CFG3 #( .INIT(8'h08) )  DataO_10_iv_0_a3_0_2 (.A(CCA_NIRQ_c), .B(
        \State2[0]_net_1 ), .C(\State2[1]_net_1 ), .Y(
        DataO_10_iv_0_a3_0_net_1));
    CFG4 #( .INIT(16'h7FFF) )  un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_x (.A(
        un1_DataI_0_a3_a_a_a_a_a_a_0_41), .B(
        un1_DataI_0_a3_a_a_a_a_a_a_0_42), .C(\Shift_reg[54]_net_1 ), 
        .D(un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_x_RNO_net_1), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_x_net_1));
    CFG4 #( .INIT(16'h8000) )  un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_RNO (
        .A(\Shift_reg[42]_net_1 ), .B(\Shift_reg[47]_net_1 ), .C(
        \Shift_reg[54]_net_1 ), .D(\Shift_reg[48]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_40));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_58_838_i_m4_ns (.A(
        Shift_reg_68_58_838_i_m4_am_net_1), .B(
        Shift_reg_68_58_838_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3511));
    SLE \TC_Error_Counter[5]  (.D(\TC_Error_Counter_s[5] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[5]));
    SLE \Shift_reg[48]  (.D(N_4627_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[48]_net_1 ));
    CFG4 #( .INIT(16'h9009) )  Shift_reg_68_46_1115_i_i_N_4L7 (.A(
        \Parity[5]_net_1 ), .B(\Syn_reg[5]_net_1 ), .C(
        \Syn_reg[6]_net_1 ), .D(\Parity[6]_net_1 ), .Y(
        Shift_reg_68_46_1115_i_i_N_4L7_net_1));
    CFG4 #( .INIT(16'h2814) )  Shift_reg_68_sn_m23_0_a2 (.A(
        \Syn_reg[5]_net_1 ), .B(\Syn_reg[2]_net_1 ), .C(
        \Parity[2]_net_1 ), .D(\Parity[5]_net_1 ), .Y(
        Shift_reg_68_sn_N_24));
    CFG4 #( .INIT(16'hFF7F) )  un1_DataI_0_a3_a_a_a_a_a_a_N_4L5 (.A(
        un1_DataI_0_a3_a_a_a_a_a_a_0_41), .B(
        un1_DataI_0_a3_a_a_a_a_a_a_0_42), .C(
        un1_DataI_0_a3_a_a_a_a_a_a_0_40), .D(
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_sx_net_1), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_N_4L5_net_1));
    CFG2 #( .INIT(4'h2) )  Start_Buff_10_7_336_a2 (.A(N_2131_1), .B(
        \State1[0]_net_1 ), .Y(N_3082));
    SLE \Parity[4]  (.D(N_3147_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_10_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Parity[4]_net_1 ));
    SLE \TC_Packet_Counter[8]  (.D(\TC_Packet_Counter_s[8] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[8]));
    CFG4 #( .INIT(16'hF5F7) )  Shift_reg_68_56_895_i_1 (.A(CCA_NIRQ_c), 
        .B(\Shift_reg[5]_net_1 ), .C(N_3562), .D(
        Shift_reg_68_sn_N_84_mux), .Y(Shift_reg_68_56_895_i_1_net_1));
    CFG4 #( .INIT(16'h3337) )  Shift_reg_68_7_2129_i_0 (.A(
        \Shift_reg[50]_net_1 ), .B(CCA_NIRQ_c), .C(
        Shift_reg_68_sn_N_56), .D(N_82), .Y(
        Shift_reg_68_7_2129_i_0_net_1));
    CFG2 #( .INIT(4'h1) )  Shift_reg_68_28_10_0_a2 (.A(
        \Bit_Counter[2]_net_1 ), .B(\Bit_Counter[1]_net_1 ), .Y(
        Shift_reg_68_28_9_2));
    SLE \TC_Error_Counter[7]  (.D(\TC_Error_Counter_s[7] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[7]));
    CFG2 #( .INIT(4'h7) )  Shift_reg_68_30_1493_i_i_o3_1_0 (.A(N_82), 
        .B(Shift_m5_0), .Y(Shift_reg_68_30_1493_i_i_o3_1_net_1));
    CFG4 #( .INIT(16'h0C84) )  Shift_reg_68_20_1753_i_a7_1_0 (.A(
        Shift_reg_68_50_9), .B(Shift_reg_68_sn_N_56), .C(
        \Shift_reg[35]_net_1 ), .D(\un1_Syn_reg[0] ), .Y(
        Shift_reg_68_20_1753_i_a7_1_0_net_1));
    CFG4 #( .INIT(16'hF780) )  Shift_reg_68_18_1811_i_m4_bm (.A(
        Shift_reg_68_28_15_0_net_1), .B(Shift_reg_68_28_41_4), .C(
        RX_GPIO0_c), .D(\Shift_reg[33]_net_1 ), .Y(
        Shift_reg_68_18_1811_i_m4_bm_net_1));
    SLE \Bit_Counter[1]  (.D(\Bit_Counter_lm[1] ), .CLK(RX_GPIO1_c), 
        .EN(un1_DataO41_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Bit_Counter[1]_net_1 ));
    CFG4 #( .INIT(16'hF0F1) )  \State1_ns_0_o5_3_RNIMTT5B[0]  (.A(
        un1_TC_Packet_Counter17_3_net_1), .B(
        \State1_ns_0_o5_2[0]_net_1 ), .C(Shift_m3_0_sx), .D(
        \State1_ns_0_o5_3[0]_net_1 ), .Y(Shift_N_5));
    CFG3 #( .INIT(8'hD8) )  Shift_reg_68_24_1637_i_0_o2_2 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_50_5), .C(N_82), .Y(
        N_272));
    CFG4 #( .INIT(16'h0015) )  \Shift_reg_RNO_1[3]  (.A(N_3606), .B(
        un1_TC_Packet_Counter17_5_net_1), .C(\State1[0]_net_1 ), .D(
        Shift_reg_68_53_953_i_0_net_1), .Y(N_3605_i_1));
    CFG4 #( .INIT(16'h10C0) )  \un1_Syn_reg_i_o3_RNIFELN_0[2]  (.A(
        \un1_Syn_reg[2] ), .B(N_53_i), .C(\un1_Syn_reg[0] ), .D(
        \un1_Syn_reg[6] ), .Y(\Shift_reg_68_54_e_0[11] ));
    SLE \TC_Error_Counter[15]  (.D(\TC_Error_Counter_s[15] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[15]));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_35_1349_i_a7_2 (.A(
        Shift_reg_68_sn_N_56), .B(\Shift_reg[19]_net_1 ), .C(N_82), .Y(
        N_3939));
    CFG4 #( .INIT(16'h084C) )  un1_Syn_reg_67_1_x2_2_i_o3_RNIVE0N3 (.A(
        \un1_Syn_reg[0] ), .B(\State1[0]_net_1 ), .C(N_2176), .D(
        Shift_reg_68_sn_N_42), .Y(Shift_reg_68_sn_N_49));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIOQSJ6[18]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[18]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[17] ), .S(
        \TC_Packet_Counter_s[18] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[18] ));
    CFG3 #( .INIT(8'h54) )  \un1_Syn_reg_i_o3_0_x2_RNIJI7CA[1]  (.A(
        Shift_reg_68_sn_m72_7_ns_sx_0), .B(N_53_i), .C(N_2548), .Y(
        Shift_reg_68_sn_N_73));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[23]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[23]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[22]_net_1 ), .S(
        \TC_Error_Counter_s[23] ), .Y(), .FCO(
        \TC_Error_Counter_cry[23]_net_1 ));
    CFG4 #( .INIT(16'h0C84) )  Shift_reg_68_11_2010_i_a7_1_0 (.A(
        Shift_reg_68_50_5), .B(Shift_reg_68_sn_N_56), .C(
        \Shift_reg[54]_net_1 ), .D(\un1_Syn_reg[0] ), .Y(
        Shift_reg_68_11_2010_i_a7_1_0_net_1));
    CFG2 #( .INIT(4'h1) )  Shift_reg_68_54 (.A(Shift_reg_68_sn_N_49), 
        .B(Shift_reg_68_sn_N_33), .Y(Shift_reg_68_54_net_1));
    CFG4 #( .INIT(16'hFFF4) )  Shift_reg_68_23_1667_i_i (.A(N_216), .B(
        N_253), .C(N_171), .D(N_172), .Y(N_63));
    SLE \Start_Buff[14]  (.D(N_3356), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[14]_net_1 ));
    SLE \Start_Buff[3]  (.D(Start_Buff_10_5_358_a2_net_1), .CLK(
        RX_GPIO1_c), .EN(un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[3]_net_1 ));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[43]  (.A(
        Shift_reg_68_28_25_0_net_1), .B(N_92), .C(RX_GPIO0_c), .D(
        \Shift_reg[43]_net_1 ), .Y(N_113));
    CFG4 #( .INIT(16'h02CC) )  \un1_Syn_reg_RNIRK8I_0[3]  (.A(
        \un1_Syn_reg[3]_net_1 ), .B(\un1_Syn_reg[2] ), .C(N_53_i), .D(
        \un1_Syn_reg[6] ), .Y(Shift_reg_68_sn_m47_0_ns_1));
    CFG4 #( .INIT(16'h50D0) )  Shift_reg_68_24_1637_i_0_0 (.A(N_62), 
        .B(N_82), .C(Shift_reg_68_24_1637_i_0_0_N_2L1_net_1), .D(
        Shift_reg_68_sn_N_56), .Y(Shift_reg_68_24_1637_i_0_0_net_1));
    CFG4 #( .INIT(16'hFFBF) )  Shift_reg_68_13_1953_i_i_o2 (.A(
        \Bit_Counter[2]_net_1 ), .B(un14lto0), .C(\State1[0]_net_1 ), 
        .D(N_58), .Y(N_87));
    CFG3 #( .INIT(8'hB3) )  Shift_reg_1_sqmuxa_1_i_o3_0_o2 (.A(N_436_1)
        , .B(TC_Packet_Counter17_i_0), .C(un14lto5), .Y(N_58));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_52_983_i_m4_ns (.A(
        Shift_reg_68_52_983_i_m4_am_net_1), .B(
        Shift_reg_68_52_983_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3630));
    SLE \Shift_reg[34]  (.D(N_4292_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[34]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \State1_ns_0_1[0]  (.A(
        \State1_ns_0_a5_2_9[0]_net_1 ), .B(Bit_Counter_3_sqmuxa), .C(
        N_2130), .D(\State1_ns_0_a5_2_8[0]_net_1 ), .Y(
        \State1_ns_0_1[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \Shift_reg_RNIS8J6[26]  (.A(
        \Shift_reg[31]_net_1 ), .B(\Shift_reg[38]_net_1 ), .C(
        \Shift_reg[32]_net_1 ), .D(\Shift_reg[26]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_38));
    CFG4 #( .INIT(16'hF5F7) )  Shift_reg_68_35_1349_i_1 (.A(CCA_NIRQ_c)
        , .B(\Shift_reg[19]_net_1 ), .C(N_3939), .D(
        Shift_reg_68_sn_N_84_mux), .Y(Shift_reg_68_35_1349_i_1_net_1));
    CFG4 #( .INIT(16'hFCEC) )  un1_DataO41_24_i_0 (.A(
        un1_DataO41_24_i_a3_0_4_net_1), .B(N_357), .C(N_295), .D(
        un1_DataO41_18_1_0_RNIGFRM_Y), .Y(N_88));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_20_1753_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_82), 
        .D(N_105), .Y(N_4275));
    CFG4 #( .INIT(16'h0F0B) )  un1_Start_Buff_1_RNIJQRQ (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(un1_CCA_i_0), .D(
        un1_Start_Buff_1_net_1), .Y(un1_DataO41_5_i_0));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_62_726_i_m4_ns (.A(
        Shift_reg_68_62_726_i_m4_am_net_1), .B(
        Shift_reg_68_62_726_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3411));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[8]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3486), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3483_i_0));
    SLE IP_END (.D(N_3002), .CLK(RX_GPIO1_c), .EN(un1_DataO41_19_i_0), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_IP_END));
    CFG4 #( .INIT(16'h6F4C) )  \Shift_reg_RNO_0[43]  (.A(
        \Shift_reg_RNO_2[43]_net_1 ), .B(\Shift_reg[43]_net_1 ), .C(
        N_349_1), .D(Shift_reg_68_sn_N_84_mux), .Y(N_4752_i_1));
    CFG4 #( .INIT(16'h0008) )  Shift_reg_68_28_47 (.A(un14lto4), .B(
        Shift_reg_68_28_9_2), .C(N_389), .D(N_57), .Y(
        Shift_reg_68_28_47_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIL8457[21]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[21]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[20] ), .S(
        \TC_Packet_Counter_s[21] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[21] ));
    CFG4 #( .INIT(16'hFE04) )  Parity_16_3_456_i_m5 (.A(
        \Parity_Counter[0]_net_1 ), .B(RX_GPIO0_c), .C(
        Parity_16_3_456_i_o4_0), .D(\Parity[2]_net_1 ), .Y(N_3190));
    CFG4 #( .INIT(16'h2000) )  \State1_ns_0_a5_2_8[0]  (.A(
        \Start_Buff[9]_net_1 ), .B(\Start_Buff[10]_net_1 ), .C(
        un1_Start_Buff_1_11_net_1), .D(un1_Start_Buff_1_5_net_1), .Y(
        \State1_ns_0_a5_2_8[0]_net_1 ));
    CFG4 #( .INIT(16'h5030) )  \un1_Syn_reg_i_o3_0_x2_RNI64E57_1[1]  (
        .A(Shift_reg_68_sn_m59_i_x3_RNI3Q7P3_net_1), .B(
        Shift_reg_68_sn_m72_6_ns_1), .C(N_53_i), .D(\un1_Syn_reg[6] ), 
        .Y(Shift_reg_68_sn_m72_7_ns_sx_0));
    CFG4 #( .INIT(16'h0040) )  un1_DataI_0_a3_a_a_a_a_a_a_x_RNO (.A(
        \Shift_reg[53]_net_1 ), .B(\Parity[4]_net_1 ), .C(
        \Parity[2]_net_1 ), .D(\Shift_reg[51]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_33));
    CFG3 #( .INIT(8'h6C) )  \Shift_reg_RNO_0[3]  (.A(Shift_reg_68_50_2)
        , .B(\Shift_reg[3]_net_1 ), .C(\un1_Syn_reg[2] ), .Y(
        N_1426_mux));
    CFG4 #( .INIT(16'h159D) )  DataO_10_iv_0_0_RNO_29 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[23]_net_1 ), .D(\Shift_reg[19]_net_1 ), .Y(
        DataO_6_3_i_m2_1_2));
    CFG4 #( .INIT(16'h0307) )  Shift_reg_68_30_1493_i_i_o3 (.A(
        Shift_reg_68_1_2300_i_0_o2), .B(
        Shift_reg_68_30_1493_i_i_o3_1_net_1), .C(Shift_N_7_mux_2), .D(
        un1_TC_Packet_Counter17_3_RNIS3QPC_net_1), .Y(N_114));
    CFG2 #( .INIT(4'h6) )  Shift_reg_68_sn_m57_i_o3 (.A(
        \Parity[5]_net_1 ), .B(\Syn_reg[5]_net_1 ), .Y(
        \un1_Syn_reg[5] ));
    SLE \Start_Buff[7]  (.D(N_3062), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[7]_net_1 ));
    SLE \Start_Buff[15]  (.D(N_3346), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[15]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  Shift_reg_68_26_1580_i_i_N_2L1 (.A(
        un14lto4), .B(\Bit_Counter[2]_net_1 ), .C(un14lto5), .D(
        un14lto0), .Y(Shift_reg_68_26_1580_i_i_N_2L1_net_1));
    CFG4 #( .INIT(16'hF66F) )  Shift_reg_68_44_0_o3 (.A(
        \Parity[5]_net_1 ), .B(\Syn_reg[5]_net_1 ), .C(
        \Syn_reg[6]_net_1 ), .D(\Parity[6]_net_1 ), .Y(N_109));
    SLE \State2[1]  (.D(State2_2_sqmuxa), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_12_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \State2[1]_net_1 ));
    CFG4 #( .INIT(16'h195D) )  DataO_10_iv_0_0_RNO_30 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[17]_net_1 ), .D(\Shift_reg[21]_net_1 ), .Y(
        DataO_6_6_i_m2_1_2));
    CFG4 #( .INIT(16'hFB40) )  Shift_reg_68_42_1143_i_m4_bm (.A(N_110), 
        .B(Shift_reg_68_28_50_4), .C(RX_GPIO0_c), .D(
        \Shift_reg[26]_net_1 ), .Y(Shift_reg_68_42_1143_i_m4_bm_net_1));
    CFG4 #( .INIT(16'h78F0) )  Shift_reg_68_2_2272_i_m4_am (.A(
        \Shift_reg_68_54_e_0[7] ), .B(Shift_reg_68_54_4), .C(
        \Shift_reg[45]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_2_2272_i_m4_am_net_1));
    CFG4 #( .INIT(16'h666F) )  Shift_reg_68_44_4_0_o3 (.A(
        \Syn_reg[6]_net_1 ), .B(\Parity[6]_net_1 ), .C(
        \un1_Syn_reg[2] ), .D(\un1_Syn_reg[3]_net_1 ), .Y(N_204));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_4_369_a2 (.A(CCA_NIRQ_c), .B(
        \Start_Buff[1]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3112));
    CFG4 #( .INIT(16'h0001) )  \Shift_reg_RNI6NN6[37]  (.A(
        \Shift_reg[44]_net_1 ), .B(\Shift_reg[49]_net_1 ), .C(
        \Shift_reg[43]_net_1 ), .D(\Shift_reg[37]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_45));
    SLE \TC_Error_Counter[2]  (.D(\TC_Error_Counter_s[2] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[2]));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[28]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[28]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[27]_net_1 ), .S(
        \TC_Error_Counter_s[28] ), .Y(), .FCO(
        \TC_Error_Counter_cry[28]_net_1 ));
    CFG2 #( .INIT(4'h4) )  State2_2_sqmuxa_0_a3 (.A(N_302), .B(
        DataO_10_iv_0_a3_0_net_1), .Y(State2_2_sqmuxa));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_8_2099_i_0_a3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_82), 
        .D(N_121), .Y(N_346));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[33]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4320), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4317_i_0));
    SLE \TC_Error_Counter[20]  (.D(\TC_Error_Counter_s[20] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[20]));
    CFG3 #( .INIT(8'hF1) )  Block_ErrO_0_sqmuxa_i_o3 (.A(
        \State1_ns_0_o5_3[0]_net_1 ), .B(\State1_ns_0_o5_2[0]_net_1 ), 
        .C(un1_TC_Packet_Counter17_3_net_1), .Y(N_295));
    CFG2 #( .INIT(4'h6) )  \un1_Syn_reg_i_o3_0_x2[1]  (.A(
        \Parity[1]_net_1 ), .B(\Syn_reg[1]_net_1 ), .Y(N_53_i));
    CFG3 #( .INIT(8'hA9) )  Shift_reg_68_47_1039_i_m4_0_am (.A(
        \Shift_reg[0]_net_1 ), .B(\un1_Syn_reg[2] ), .C(N_204), .Y(
        Shift_reg_68_47_1039_i_m4_0_am_net_1));
    CFG3 #( .INIT(8'hBF) )  Shift_reg_68_37_1293_i_0_o3 (.A(
        Shift_reg_68_37_1293_i_0_o3_1_net_1), .B(
        \Bit_Counter[1]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_402));
    CFG4 #( .INIT(16'hAAFE) )  un1_DataO41_18_1_RNI2TCP (.A(
        un1_DataO41_18_1_net_1), .B(\State1_ns_0_o5_3[0]_net_1 ), .C(
        \State1_ns_0_o5_2[0]_net_1 ), .D(
        un1_TC_Packet_Counter17_3_net_1), .Y(un1_DataO41_18));
    ARI1 #( .INIT(20'h4AA00) )  TC_Error_Counter_s_367 (.A(VCC_net_1), 
        .B(CLTU_0_TC_Error_Counter[0]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(VCC_net_1), .S(), .Y(), .FCO(TC_Error_Counter_s_367_FCO));
    CFG4 #( .INIT(16'h37F7) )  Shift_reg_68_30_1493_i_i_0_RNO (.A(
        N_122), .B(\Shift_reg[14]_net_1 ), .C(N_82), .D(N_210), .Y(
        Shift_N_9_0));
    SLE \Shift_Bit_Counter[2]  (.D(\Shift_Bit_Counter_s[2] ), .CLK(
        RX_GPIO1_c), .EN(Shift_Bit_Countere), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \un22_DataO_i[2] ));
    CFG4 #( .INIT(16'h7362) )  DataO_10_iv_0_a3_0_RNO_6 (.A(
        \un6_DataO_i[3] ), .B(DataO_2_3_1_2), .C(
        \Start_Buff[15]_net_1 ), .D(\Start_Buff[11]_net_1 ), .Y(N_2617)
        );
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h0080) )  Shift_reg_68_28_13 (.A(
        \Bit_Counter[3]_net_1 ), .B(Shift_reg_68_28_17_2), .C(
        Shift_reg_68_28_9_2), .D(N_57), .Y(Shift_reg_68_28_13_net_1));
    CFG4 #( .INIT(16'h2000) )  \un1_Syn_reg_i_o3_RNIFELN[2]  (.A(
        \un1_Syn_reg[2] ), .B(N_53_i), .C(\un1_Syn_reg[0] ), .D(
        \un1_Syn_reg[6] ), .Y(\Shift_reg_68_54_e_0[42] ));
    CFG4 #( .INIT(16'h3323) )  Shift_reg_68_9_2070_i_0_a3 (.A(
        Shift_reg_68_sn_N_56), .B(\Shift_reg[52]_net_1 ), .C(
        Shift_reg_68_sn_N_84_mux), .D(N_81), .Y(N_283));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[50]  (.A(
        Shift_reg_68_28_5_1_net_1), .B(N_86), .C(RX_GPIO0_c), .D(
        \Shift_reg[50]_net_1 ), .Y(N_120));
    CFG4 #( .INIT(16'hFCF5) )  Shift_reg_68_7_2129_i_2 (.A(
        \Shift_reg[50]_net_1 ), .B(Shift_reg_68_7_2129_i_a7_1_0_net_1), 
        .C(Shift_reg_68_7_2129_i_0_net_1), .D(Shift_reg_68_sn_N_84_mux)
        , .Y(Shift_reg_68_7_2129_i_2_net_1));
    SLE \TC_Error_Counter[16]  (.D(\TC_Error_Counter_s[16] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[16]));
    CFG4 #( .INIT(16'h0F53) )  DataO_6_53_am_1_1 (.A(
        \Shift_reg[27]_net_1 ), .B(\Shift_reg[31]_net_1 ), .C(
        \un22_DataO_i[2] ), .D(\un22_DataO_i[1] ), .Y(
        DataO_6_53_am_1_1_net_1));
    SLE \TC_Error_Counter[11]  (.D(\TC_Error_Counter_s[11] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[11]));
    CFG4 #( .INIT(16'hFFFB) )  Shift_reg_68_60_782_i_i_o2_1 (.A(
        un14lto0), .B(\Bit_Counter[2]_net_1 ), .C(N_57), .D(N_103), .Y(
        N_220));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIJU4S7[25]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[25]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[24] ), .S(
        \TC_Packet_Counter_s[25] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[25] ));
    SLE \Shift_reg[35]  (.D(N_4270_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[35]_net_1 ));
    CFG3 #( .INIT(8'h02) )  Shift_reg_68_28_31_0 (.A(
        Shift_reg_68_28_30_3), .B(N_389), .C(un14lto4), .Y(
        Shift_reg_68_28_31_0_net_1));
    CFG4 #( .INIT(16'h6030) )  Shift_reg_68_10_2040_i_a7_1 (.A(N_53_i), 
        .B(\Shift_reg[53]_net_1 ), .C(N_349_1), .D(N_1463), .Y(N_4514));
    CFG3 #( .INIT(8'hD5) )  Syn_reg_23_639_i_0_o3 (.A(CCA_NIRQ_c), .B(
        \State1[0]_net_1 ), .C(TC_Packet_Counter18_i_0), .Y(N_54));
    CFG4 #( .INIT(16'h4657) )  DataO_10_iv_0_a3_0_RNO_2 (.A(
        \un6_DataO_i[1] ), .B(\un6_DataO_i[0] ), .C(N_2620), .D(N_2617)
        , .Y(DataO_2_15_1_2));
    SLE \Start_Buff[8]  (.D(N_3052), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[8]_net_1 ));
    SLE \Start_Buff[10]  (.D(N_3032), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[10]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  Shift_reg_68_24_1637_i_0_2 (.A(
        Shift_reg_68_24_1637_i_0_a3_1_0_net_1), .B(
        Shift_reg_68_24_1637_i_0_0_net_1), .C(N_74), .D(
        Shift_reg_68_sn_N_84_mux), .Y(Shift_reg_68_24_1637_i_0_2_net_1)
        );
    CFG4 #( .INIT(16'h0AFC) )  DataO_10_iv_0_0_RNO_8 (.A(
        \Shift_reg[45]_net_1 ), .B(\Shift_reg[41]_net_1 ), .C(
        \Shift_Bit_Counter[5]_net_1 ), .D(DataO_6_37_i_m2_1_2), .Y(
        N_318));
    SLE \Start_Buff[4]  (.D(N_3092), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[4]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNI5FBI1[1]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[1]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Packet_Counter_cry[0] ), .S(
        \TC_Packet_Counter_s[1] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[1] ));
    SLE \TC_Packet_Counter[17]  (.D(\TC_Packet_Counter_s[17] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[17]));
    CFG4 #( .INIT(16'h159D) )  DataO_10_iv_0_0_RNO_22 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[4]_net_1 ), .D(\Shift_reg[0]_net_1 ), .Y(
        DataO_6_29_i_m2_0_5));
    CFG4 #( .INIT(16'hFB40) )  Shift_reg_68_52_983_i_m4_bm (.A(N_102), 
        .B(Shift_reg_68_28_42_4), .C(RX_GPIO0_c), .D(
        \Shift_reg[2]_net_1 ), .Y(Shift_reg_68_52_983_i_m4_bm_net_1));
    SLE \Shift_reg[0]  (.D(N_3677_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[0]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \Shift_reg_RNIEM0F[16]  (.A(
        \Shift_reg[16]_net_1 ), .B(\Shift_reg[18]_net_1 ), .C(
        \Shift_reg[15]_net_1 ), .D(\Shift_reg[8]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_36));
    CFG4 #( .INIT(16'h00C8) )  un1_TC_Packet_Counter17_3_RNIS3QPC (.A(
        un1_TC_Packet_Counter17_3_net_1), .B(\State1[0]_net_1 ), .C(
        Shift_m6_i_a4_1), .D(Shift_reg_68_sn_N_56), .Y(
        un1_TC_Packet_Counter17_3_RNIS3QPC_net_1));
    CFG4 #( .INIT(16'h0800) )  Shift_reg_68_28_36 (.A(
        \Bit_Counter[2]_net_1 ), .B(\Bit_Counter[1]_net_1 ), .C(N_86), 
        .D(N_436_1), .Y(Shift_reg_68_28_36_net_1));
    CFG4 #( .INIT(16'h89FF) )  Shift_reg_68_1_2300_i_0_o3_0_0 (.A(
        \un1_Syn_reg[0] ), .B(\un1_Syn_reg[6] ), .C(
        Shift_reg_68_sn_N_24), .D(N_53_i), .Y(
        Shift_reg_68_1_2300_i_0_o3_0_0_net_1));
    CFG4 #( .INIT(16'h8000) )  un1_Start_Buff_1 (.A(
        un1_Start_Buff_1_4_net_1), .B(un1_Start_Buff_1_6_net_1), .C(
        un1_Start_Buff_1_5_0), .D(un1_Start_Buff_1_11_net_1), .Y(
        un1_Start_Buff_1_net_1));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_9_2070_i_0_a3_1 (.A(N_86), .B(
        RX_GPIO0_c), .C(Shift_reg_68_9_2070_i_0_o2_1_1_net_1), .Y(
        N_286));
    CFG4 #( .INIT(16'h7362) )  DataO_10_iv_0_a3_0_RNO_0 (.A(
        \un6_DataO_i[3] ), .B(DataO_2_13_1_2), .C(
        \Start_Buff[12]_net_1 ), .D(\Start_Buff[8]_net_1 ), .Y(N_2627));
    CFG3 #( .INIT(8'h20) )  Shift_reg_68_28_17_0 (.A(
        Shift_reg_68_28_30_3), .B(un14lto5), .C(Shift_reg_68_28_17_2), 
        .Y(Shift_reg_68_28_17_0_net_1));
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_14_1925_i_m4_bm (.A(
        Shift_reg_68_28_11_0_net_1), .B(N_374), .C(RX_GPIO0_c), .D(
        \Shift_reg[29]_net_1 ), .Y(Shift_reg_68_14_1925_i_m4_bm_net_1));
    CFG3 #( .INIT(8'hFB) )  Shift_reg_68_37_1293_i_0_o3_1 (.A(N_389), 
        .B(TC_Packet_Counter17_i_0), .C(N_387), .Y(
        Shift_reg_68_37_1293_i_0_o3_1_net_1));
    CFG4 #( .INIT(16'h0400) )  Shift_reg_68_11_2010_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_124), 
        .D(N_82), .Y(N_4494));
    CFG4 #( .INIT(16'hF780) )  \Shift_reg_5[25]  (.A(
        un39_Shift_reg_0_net_1), .B(N_436_1), .C(RX_GPIO0_c), .D(
        \Shift_reg[25]_net_1 ), .Y(\Shift_reg_5[25]_net_1 ));
    SLE \TC_Packet_Counter[26]  (.D(\TC_Packet_Counter_s[26] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[26]));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[53]  (.A(
        Shift_reg_68_28_8_0_net_1), .B(N_374), .C(RX_GPIO0_c), .D(
        \Shift_reg[53]_net_1 ), .Y(N_123_0));
    CFG4 #( .INIT(16'h0007) )  \Shift_reg_RNO[54]  (.A(
        \State1[0]_net_1 ), .B(un1_TC_Packet_Counter17_5_net_1), .C(
        N_4494), .D(Shift_reg_68_11_2010_i_2_net_1), .Y(N_4489_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNI1NC05[9]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[9]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Packet_Counter_cry[8] ), .S(
        \TC_Packet_Counter_s[9] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[9] ));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[18]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3960), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3957_i_0));
    SLE \TC_Error_Counter[28]  (.D(\TC_Error_Counter_s[28] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[28]));
    CFG2 #( .INIT(4'h8) )  \block_counter_RNIKA3D[0]  (.A(
        \un1_block_counter_4[0]_net_1 ), .B(\block_counter[0]_net_1 ), 
        .Y(CO0));
    SLE \TC_Packet_Counter[21]  (.D(\TC_Packet_Counter_s[21] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[21]));
    CFG4 #( .INIT(16'hFFFE) )  Shift_reg_68_26_1580_i_i_o3 (.A(
        un14lto0), .B(N_92), .C(un14lto4), .D(un14lto5), .Y(N_219));
    CFG2 #( .INIT(4'hE) )  Shift_reg_68_1_2300_i_0_o3_1_0 (.A(N_385), 
        .B(N_91), .Y(Shift_reg_68_1_2300_i_0_o3_1_0_net_1));
    CFG2 #( .INIT(4'h8) )  TC_Packet_Counter18_i_a3_0 (.A(un14lto5), 
        .B(un14lto4), .Y(N_21_i));
    SLE \Start_Buff[11]  (.D(N_3022), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_26_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[11]_net_1 ));
    CFG3 #( .INIT(8'h20) )  Shift_reg_68_28_16 (.A(
        Shift_reg_68_28_42_4), .B(un14lto5), .C(Shift_reg_68_28_30_3), 
        .Y(Shift_reg_68_28_16_net_1));
    CFG3 #( .INIT(8'h13) )  \Shift_reg_RNO[25]  (.A(
        un1_TC_Packet_Counter17_5_net_1), .B(
        Shift_reg_68_41_1171_i_3_net_1), .C(\State1[0]_net_1 ), .Y(
        N_3792_i_0));
    CFG3 #( .INIT(8'h10) )  Shift_reg_68_26_1580_i_i_N_6L11_RNO_0 (.A(
        Shift_reg_68_1_2300_i_0_o2), .B(\Shift_reg[41]_net_1 ), .C(
        N_53_i), .Y(Shift_m3_2_1));
    CFG4 #( .INIT(16'h4800) )  un1_DataO41_22_0_a2 (.A(
        \un1_Syn_reg[2] ), .B(N_94_i), .C(\un1_Syn_reg[4] ), .D(
        \un1_Syn_reg[3]_net_1 ), .Y(N_372));
    CFG4 #( .INIT(16'h3230) )  \Shift_reg_RNO[39]  (.A(
        Shift_reg_68_sn_N_84_mux), .B(Shift_reg_68_24_1637_i_0_2_net_1)
        , .C(\Shift_reg[39]_net_1 ), .D(N_272), .Y(N_4176_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[2]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[2]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[1]_net_1 ), .S(
        \TC_Error_Counter_s[2] ), .Y(), .FCO(
        \TC_Error_Counter_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNILPHH5[12]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[12]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[11] ), .S(
        \TC_Packet_Counter_s[12] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[12] ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[21]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[21]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[20]_net_1 ), .S(
        \TC_Error_Counter_s[21] ), .Y(), .FCO(
        \TC_Error_Counter_cry[21]_net_1 ));
    CFG4 #( .INIT(16'h153F) )  \Shift_reg_RNO_1[43]  (.A(
        \Shift_reg_RNO_3[43]_net_1 ), .B(\State1[0]_net_1 ), .C(
        un1_TC_Packet_Counter17_5_net_1), .D(Shift_reg_68_sn_N_84_mux), 
        .Y(\Shift_reg_RNO_1[43]_net_1 ));
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_22_1695_i_m4_bm (.A(
        Shift_reg_68_28_19_0_net_1), .B(N_374), .C(RX_GPIO0_c), .D(
        \Shift_reg[37]_net_1 ), .Y(Shift_reg_68_22_1695_i_m4_bm_net_1));
    CFG4 #( .INIT(16'h00DC) )  Shift_reg_68_13_1953_i_i_o3_0_0 (.A(
        \un1_Syn_reg[0] ), .B(N_91), .C(N_57), .D(
        Shift_reg_68_1_2300_i_0_o2), .Y(
        Shift_reg_68_13_1953_i_i_o3_0_0_0));
    CFG3 #( .INIT(8'h47) )  \un1_Syn_reg_i_o3_0_x2_RNIAUM3A[1]  (.A(
        N_2551), .B(N_53_i), .C(N_2548), .Y(Shift_m6_i_a4_1));
    CFG4 #( .INIT(16'hFBFF) )  Shift_reg_68_13_1953_i_i_o3 (.A(
        \Bit_Counter[2]_net_1 ), .B(un14lto4), .C(N_57), .D(un14lto0), 
        .Y(N_90));
    SLE \TC_Error_Counter[27]  (.D(\TC_Error_Counter_s[27] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[27]));
    SLE \Shift_reg[50]  (.D(N_4580_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[50]_net_1 ));
    CFG2 #( .INIT(4'h8) )  Shift_reg_68_28_32_2 (.A(un14lto5), .B(
        \Bit_Counter[1]_net_1 ), .Y(Shift_reg_68_28_32_2_net_1));
    SLE \Shift_Bit_Counter[3]  (.D(\Shift_Bit_Counter_s[3] ), .CLK(
        RX_GPIO1_c), .EN(Shift_Bit_Countere), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_Bit_Counter[3]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  un1_DataO41_24_i_a3_0_1_0 (.A(
        \un6_DataO_i[0] ), .B(\un6_DataO_i[1] ), .C(\un6_DataO_i[3] ), 
        .D(\un6_DataO_i[2] ), .Y(un1_DataO41_24_i_a3_0_1_net_1));
    CFG3 #( .INIT(8'h13) )  DataO_RNO (.A(DataO_0_sqmuxa_1_0_net_1), 
        .B(un1_CCA_i_0), .C(un1_State1_1_net_1), .Y(un1_DataO41_14_i_0)
        );
    CFG4 #( .INIT(16'h0A08) )  \State2_RNO[0]  (.A(
        State2_1_sqmuxa_net_1), .B(\State1_ns_0_o5_2[0]_net_1 ), .C(
        un1_TC_Packet_Counter17_3_net_1), .D(
        \State1_ns_0_o5_3[0]_net_1 ), .Y(\State2_9[0] ));
    CFG4 #( .INIT(16'h5551) )  Shift_reg_68_63_697_i_i_N_5L8_RNO (.A(
        Shift_reg_68_1_2300_i_0_o2), .B(\State1[0]_net_1 ), .C(
        un1_TC_Packet_Counter17_3_net_1), .D(
        \State1_ns_0_o5_2[0]_net_1 ), .Y(Shift_m8_i_a3_0_sx));
    CFG2 #( .INIT(4'h7) )  Shift_reg_68_28_26_2_i (.A(un14lto5), .B(
        \Bit_Counter[3]_net_1 ), .Y(N_34));
    CFG3 #( .INIT(8'h0E) )  \un1_Start_Sequence_counter_1.SUM_m2_e  (
        .A(\State1_ns_0_o5_3[0]_net_1 ), .B(
        \State1_ns_0_o5_2[0]_net_1 ), .C(
        un1_TC_Packet_Counter17_3_net_1), .Y(SUM_m2_e));
    CFG4 #( .INIT(16'h8000) )  un1_Start_Buff_1_4 (.A(
        \Start_Buff[14]_net_1 ), .B(\Start_Buff[9]_net_1 ), .C(
        \Start_Buff[15]_net_1 ), .D(\Start_Buff[4]_net_1 ), .Y(
        un1_Start_Buff_1_4_net_1));
    CFG2 #( .INIT(4'h4) )  un1_Syn_reg_2_0_a3_RNI1MRK (.A(
        un1_Syn_reg_2), .B(\State1[0]_net_1 ), .Y(Shift_m3_e_0));
    CFG2 #( .INIT(4'h8) )  \Bit_Counter_lm_0[3]  (.A(
        Bit_Counter_3_sqmuxa), .B(\Bit_Counter_s[3] ), .Y(
        \Bit_Counter_lm[3] ));
    CFG3 #( .INIT(8'hFE) )  \un1_block_counter_7_am[0]  (.A(
        \block_counter[2]_net_1 ), .B(\block_counter[1]_net_1 ), .C(
        \block_counter[0]_net_1 ), .Y(
        \un1_block_counter_7_am[0]_net_1 ));
    CFG4 #( .INIT(16'h0AFC) )  DataO_10_iv_0_0_RNO_13 (.A(
        \Shift_reg[36]_net_1 ), .B(\Shift_reg[32]_net_1 ), .C(
        \Shift_Bit_Counter[5]_net_1 ), .D(DataO_6_29_i_m2_0_5), .Y(
        N_340));
    SLE \Parity[3]  (.D(N_3167_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_10_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Parity[3]_net_1 ));
    CFG4 #( .INIT(16'h6CCC) )  \Shift_reg_RNO_1[51]  (.A(N_53_i), .B(
        \Shift_reg[51]_net_1 ), .C(Shift_reg_68_50_9), .D(N_417_1), .Y(
        N_1463_mux));
    ARI1 #( .INIT(20'h4AA00) )  \Bit_Counter_s[5]  (.A(VCC_net_1), .B(
        un14lto5), .C(GND_net_1), .D(GND_net_1), .FCI(
        \Bit_Counter_cry[4]_net_1 ), .S(\Bit_Counter_s[5]_net_1 ), .Y()
        , .FCO());
    CFG4 #( .INIT(16'hF078) )  Shift_reg_68_51_1011_i_m4_am (.A(
        \Shift_reg_68_54_e_0[1] ), .B(Shift_reg_68_54_2), .C(
        \Shift_reg[1]_net_1 ), .D(\un1_Syn_reg[2] ), .Y(
        Shift_reg_68_51_1011_i_m4_am_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIOFL78[27]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[27]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[26] ), .S(
        \TC_Packet_Counter_s[27] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[27] ));
    SLE \Bit_Counter[2]  (.D(\Bit_Counter_lm[2] ), .CLK(RX_GPIO1_c), 
        .EN(un1_DataO41_5_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Bit_Counter[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  Shift_reg_68_28_19_0 (.A(N_55), .B(
        Shift_reg_68_28_17_2), .Y(Shift_reg_68_28_19_0_net_1));
    CFG4 #( .INIT(16'hF5F7) )  Shift_reg_68_17_1839_i_1 (.A(CCA_NIRQ_c)
        , .B(\Shift_reg[32]_net_1 ), .C(N_4346), .D(
        Shift_reg_68_sn_N_84_mux), .Y(Shift_reg_68_17_1839_i_1_net_1));
    SLE \Shift_reg[33]  (.D(N_4317_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[33]_net_1 ));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[20]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_3913), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_3910_i_0));
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_55_925_i_m4_bm (.A(
        Shift_reg_68_28_32_2_net_1), .B(N_90), .C(RX_GPIO0_c), .D(
        \Shift_reg[4]_net_1 ), .Y(Shift_reg_68_55_925_i_m4_bm_net_1));
    CFG4 #( .INIT(16'hF078) )  Shift_reg_68_4_2216_i_m4_am (.A(
        \Shift_reg_68_54_e_0[29] ), .B(Shift_reg_68_54_4), .C(
        \Shift_reg[47]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_4_2216_i_m4_am_net_1));
    CFG4 #( .INIT(16'h0002) )  Shift_reg_68_46_1115_i_i_N_8L17_1_RNO (
        .A(Shift_m3_e_0), .B(N_2843), .C(N_2847), .D(N_2846), .Y(
        Shift_m3_e_3));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[31]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4367), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4364_i_0));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[5]  (.A(
        Shift_reg_68_28_45_0_net_1), .B(N_374), .C(RX_GPIO0_c), .D(
        \Shift_reg[5]_net_1 ), .Y(N_75_0));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[23]  (.A(
        Shift_reg_68_28_35_1_net_1), .B(N_57), .C(RX_GPIO0_c), .D(
        \Shift_reg[23]_net_1 ), .Y(N_93));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[26]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[26]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[25]_net_1 ), .S(
        \TC_Error_Counter_s[26] ), .Y(), .FCO(
        \TC_Error_Counter_cry[26]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_15_1897_i_m4_ns (.A(
        Shift_reg_68_15_1897_i_m4_am_net_1), .B(
        Shift_reg_68_15_1897_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4392));
    CFG2 #( .INIT(4'h4) )  \Syn_reg_RNI68SL1[1]  (.A(
        Shift_reg_68_sn_N_16), .B(Shift_reg_68_sn_N_78_mux), .Y(
        \Shift_reg_68_54_e_0[17] ));
    CFG2 #( .INIT(4'h1) )  Shift_reg_68_28_16_3 (.A(
        \Bit_Counter[3]_net_1 ), .B(\Bit_Counter[1]_net_1 ), .Y(
        Shift_reg_68_28_30_3));
    CFG4 #( .INIT(16'h3337) )  Shift_reg_68_10_2040_i_0 (.A(
        \Shift_reg[53]_net_1 ), .B(CCA_NIRQ_c), .C(
        Shift_reg_68_sn_N_56), .D(N_82), .Y(N_4511_i_1_1));
    CFG4 #( .INIT(16'h195D) )  DataO_10_iv_0_0_RNO_17 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[9]_net_1 ), .D(\Shift_reg[13]_net_1 ), .Y(
        DataO_6_37_i_m2_1_2));
    CFG4 #( .INIT(16'hFF2F) )  Shift_reg_68_13_1953_i_i (.A(
        \Shift_reg[28]_net_1 ), .B(
        Shift_reg_68_1_2300_i_0_o2_0_RNIHMNKG_net_1), .C(
        Shift_reg_68_13_1953_i_i_1), .D(
        Shift_reg_68_13_1953_i_i_0_net_1), .Y(N_61));
    CFG4 #( .INIT(16'h0001) )  \Shift_reg_RNO[52]  (.A(N_285), .B(
        N_283), .C(N_286), .D(N_74), .Y(N_4533_i_0));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_31_1463_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_82), 
        .D(N_85), .Y(N_4037));
    CFG4 #( .INIT(16'h3020) )  Shift_reg_68_21_1723_i_i_a2_1_0 (.A(
        N_90), .B(Shift_reg_68_sn_N_56), .C(\Shift_reg[36]_net_1 ), .D(
        N_100), .Y(Shift_reg_68_21_1723_i_i_a2_1));
    CFG4 #( .INIT(16'hFCDC) )  un1_DataO41_27_a1_0_RNIETU41 (.A(
        \State1[0]_net_1 ), .B(un1_CCA_i_0), .C(
        Syn_reg_0_sqmuxa_2_net_1), .D(un1_DataO41_27_a1_0_net_1), .Y(
        un1_DataO41_1));
    CFG4 #( .INIT(16'hFCF5) )  Shift_reg_68_41_1171_i_3 (.A(
        \Shift_reg[25]_net_1 ), .B(Shift_reg_68_41_1171_i_a7_0_1_net_1)
        , .C(Shift_reg_68_41_1171_i_1_net_1), .D(
        Shift_reg_68_sn_N_84_mux), .Y(Shift_reg_68_41_1171_i_3_net_1));
    CFG4 #( .INIT(16'h0F22) )  Shift_reg_68_sn_m59_i_x3_RNI4RG33 (.A(
        N_54_i), .B(N_404), .C(N_41), .D(\un1_Syn_reg[0] ), .Y(
        Shift_reg_68_sn_m72_6_ns_1));
    CFG3 #( .INIT(8'h82) )  Shift_reg_68_sn_m59_i_x3_RNI590H (.A(
        N_54_i), .B(\un1_Syn_reg[2] ), .C(\un1_Syn_reg[3]_net_1 ), .Y(
        Shift_reg_68_sn_m59_i_x3_RNI590H_net_1));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_22_1695_i_m4_ns (.A(
        Shift_reg_68_22_1695_i_m4_am_net_1), .B(
        Shift_reg_68_22_1695_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4226));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_8_325_a2 (.A(CCA_NIRQ_c), .B(
        \Start_Buff[5]_net_1 ), .C(\State1[0]_net_1 ), .Y(N_3072));
    CFG4 #( .INIT(16'hFE10) )  Parity_16_5_407_i_m5 (.A(
        \Parity_Counter[0]_net_1 ), .B(Parity_16_5_407_i_o4_0_net_1), 
        .C(RX_GPIO0_c), .D(\Parity[4]_net_1 ), .Y(N_3150));
    CFG3 #( .INIT(8'hD8) )  Shift_reg_68_5_2187_i_m4_0_ns (.A(N_82), 
        .B(N_118), .C(N_206), .Y(N_4629));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_56_895_i_a7_2 (.A(
        Shift_reg_68_sn_N_56), .B(\Shift_reg[5]_net_1 ), .C(N_82), .Y(
        N_3562));
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_36_1321_i_m4_RNO_0 (.A(
        Shift_reg_68_28_32_0_net_1), .B(N_86), .C(RX_GPIO0_c), .D(
        \Shift_reg[20]_net_1 ), .Y(N_1429_mux));
    CFG2 #( .INIT(4'h6) )  \un1_Syn_reg_i_o3[2]  (.A(\Parity[2]_net_1 )
        , .B(\Syn_reg[2]_net_1 ), .Y(\un1_Syn_reg[2] ));
    CFG4 #( .INIT(16'h8000) )  \Shift_reg_RNIJTKN[10]  (.A(
        \Shift_reg[14]_net_1 ), .B(\Shift_reg[6]_net_1 ), .C(
        \Shift_reg[10]_net_1 ), .D(\Shift_reg[7]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_35));
    SLE \TC_Packet_Counter[25]  (.D(\TC_Packet_Counter_s[25] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[25]));
    CFG4 #( .INIT(16'h0080) )  Shift_reg_68_28_14_0 (.A(
        \Bit_Counter[1]_net_1 ), .B(\Bit_Counter[2]_net_1 ), .C(
        un14lto0), .D(N_57), .Y(Shift_reg_68_28_3_4));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[12]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[12]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[11]_net_1 ), .S(
        \TC_Error_Counter_s[12] ), .Y(), .FCO(
        \TC_Error_Counter_cry[12]_net_1 ));
    CFG4 #( .INIT(16'h0008) )  Shift_reg_68_sn_m57_i_o3_RNIFLIB (.A(
        \un1_Syn_reg[5] ), .B(\un1_Syn_reg[2] ), .C(\un1_Syn_reg[6] ), 
        .D(N_53_i), .Y(Shift_reg_68_sn_N_82_mux));
    CFG4 #( .INIT(16'hFFFE) )  Shift_reg_68_6_2159_i_i_o3 (.A(un14lto4)
        , .B(un14lto0), .C(N_100), .D(N_92), .Y(N_217));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[20]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[20]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[19]_net_1 ), .S(
        \TC_Error_Counter_s[20] ), .Y(), .FCO(
        \TC_Error_Counter_cry[20]_net_1 ));
    CFG4 #( .INIT(16'hF0B8) )  Shift_reg_68_47_1039_i_m4 (.A(N_3679), 
        .B(Shift_reg_68_sn_N_84_mux), .C(\Shift_reg[0]_net_1 ), .D(
        Shift_reg_68_sn_N_56), .Y(N_3680));
    SLE \block_counter[1]  (.D(\block_counter_8[1]_net_1 ), .CLK(
        RX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \block_counter[1]_net_1 ));
    CFG4 #( .INIT(16'h7030) )  Shift_reg_68_21_1723_i_i_a2_6 (.A(
        un1_TC_Packet_Counter17_3_net_1), .B(\State1[0]_net_1 ), .C(
        Shift_reg_68_21_1723_i_i_a2_6_1_net_1), .D(
        Shift_reg_68_sn_N_73), .Y(N_250));
    CFG4 #( .INIT(16'hA0DD) )  DataO_10_iv_0_0_RNO (.A(
        \Shift_Bit_Counter[3]_net_1 ), .B(N_2682), .C(N_2675), .D(
        DataO_6_55_i_m2_1_2), .Y(N_309));
    CFG3 #( .INIT(8'h04) )  \Shift_reg_RNO_3[43]  (.A(
        Shift_reg_68_sn_N_56), .B(N_82), .C(N_113), .Y(
        \Shift_reg_RNO_3[43]_net_1 ));
    SLE \Shift_reg[20]  (.D(N_3910_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[20]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \Syn_reg_RNO[4]  (.A(N_54), .B(
        \Syn_reg[3]_net_1 ), .Y(N_3275_i_0));
    SLE \TC_Error_Counter[12]  (.D(\TC_Error_Counter_s[12] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[12]));
    CFG4 #( .INIT(16'h0100) )  
        Shift_reg_68_0_2328_i_a7_0_0_a3_0_a3_0_a2_1_1 (.A(N_2846), .B(
        N_2847), .C(
        Shift_reg_68_0_2328_i_a7_0_0_a3_0_a3_0_a2_1_1_sx_net_1), .D(
        Shift_m3_e_0), .Y(
        Shift_reg_68_0_2328_i_a7_0_0_a3_0_a3_0_a2_1_1_net_1));
    CFG3 #( .INIT(8'h08) )  Start_Buff_10_3_380_a2 (.A(CCA_NIRQ_c), .B(
        \Start_Buff[0]_net_1 ), .C(\State1[0]_net_1 ), .Y(
        Start_Buff_10_3_380_a2_net_1));
    CFG2 #( .INIT(4'hB) )  Shift_reg_68_28_27_0_a2_i_o2 (.A(un14lto0), 
        .B(un14lto5), .Y(N_389));
    CFG4 #( .INIT(16'h2A3F) )  Shift_reg_68_26_1580_i_i_N_6L11 (.A(
        Shift_N_5), .B(N_253), .C(Shift_reg_68_26_1580_i_i_N_4L6_net_1)
        , .D(Shift_m3_2_3), .Y(Shift_reg_68_26_1580_i_i_1_1));
    CFG4 #( .INIT(16'hFD20) )  Shift_reg_68_15_1897_i_m4_bm (.A(
        Shift_reg_68_28_12_0_net_1), .B(N_86), .C(RX_GPIO0_c), .D(
        \Shift_reg[30]_net_1 ), .Y(Shift_reg_68_15_1897_i_m4_bm_net_1));
    CFG4 #( .INIT(16'h1115) )  un1_State1_0_RNI2E5C1 (.A(un1_CCA_i_0), 
        .B(State2_1_sqmuxa_net_1), .C(un1_State1_0_net_1), .D(
        TC_Packet_Counter19_net_1), .Y(un1_DataO41_12_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNII00T5[14]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[14]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[13] ), .S(
        \TC_Packet_Counter_s[14] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[14] ));
    CFG3 #( .INIT(8'hD8) )  Shift_reg_68_32_1435_i_m4_bm (.A(
        Shift_reg_68_28_28_net_1), .B(RX_GPIO0_c), .C(
        \Shift_reg[16]_net_1 ), .Y(Shift_reg_68_32_1435_i_m4_bm_net_1));
    CFG4 #( .INIT(16'h9669) )  \Syn_reg_RNIUMFH1_0[3]  (.A(
        \Syn_reg[3]_net_1 ), .B(\Parity[3]_net_1 ), .C(
        \Syn_reg[2]_net_1 ), .D(\Parity[2]_net_1 ), .Y(N_376));
    CFG4 #( .INIT(16'h0040) )  Shift_reg_68_53_953_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_82), 
        .D(N_73_0), .Y(N_3610));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIS6S44[7]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[7]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Packet_Counter_cry[6] ), .S(
        \TC_Packet_Counter_s[7] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[7] ));
    CFG4 #( .INIT(16'h4000) )  Shift_reg_68_6_2159_i_i_a2 (.A(N_74), 
        .B(Shift_reg_68_sn_N_84_mux), .C(\Shift_reg[49]_net_1 ), .D(
        N_217), .Y(N_231));
    SLE \TC_Error_Counter[8]  (.D(\TC_Error_Counter_s[8] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[8]));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_42_1143_i_m4_ns (.A(
        Shift_reg_68_42_1143_i_m4_am_net_1), .B(
        Shift_reg_68_42_1143_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3770));
    CFG4 #( .INIT(16'h0008) )  Shift_reg_68_28_27 (.A(
        Shift_reg_68_28_9_2), .B(\Bit_Counter[3]_net_1 ), .C(N_57), .D(
        N_389), .Y(Shift_reg_68_28_27_net_1));
    CFG4 #( .INIT(16'h7362) )  DataO_10_iv_0_a3_0_RNO_5 (.A(
        \un6_DataO_i[3] ), .B(DataO_2_6_1_2), .C(
        \Start_Buff[13]_net_1 ), .D(\Start_Buff[9]_net_1 ), .Y(N_2620));
    SLE \TC_Error_Counter[29]  (.D(\TC_Error_Counter_s[29] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[29]));
    CFG2 #( .INIT(4'h6) )  un1_Syn_reg_67_1_x2_2_i_o3 (.A(
        \Parity[0]_net_1 ), .B(\Syn_reg[0]_net_1 ), .Y(
        \un1_Syn_reg[0] ));
    CFG1 #( .INIT(2'h1) )  \TC_Error_Counter_RNO[0]  (.A(
        CLTU_0_TC_Error_Counter[0]), .Y(\TC_Error_Counter_s[0] ));
    CFG2 #( .INIT(4'h1) )  Shift_reg_68_28_15_3 (.A(un14lto0), .B(
        \Bit_Counter[3]_net_1 ), .Y(Shift_reg_68_28_29_3));
    SLE \TC_Error_Counter[3]  (.D(\TC_Error_Counter_s[3] ), .CLK(
        RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[3]));
    CFG2 #( .INIT(4'h1) )  \State1_ns_0_a5_1_0[0]  (.A(
        \block_counter[2]_net_1 ), .B(CCA_NIRQ_c), .Y(
        \State1_ns_0_a5_1_0[0]_net_1 ));
    CFG4 #( .INIT(16'h7FAF) )  Shift_reg_68_26_1580_i_i (.A(
        \Shift_reg[41]_net_1 ), .B(
        Shift_reg_68_1_2300_i_0_o2_0_RNIHMNKG_net_1), .C(
        Shift_reg_68_26_1580_i_i_1_1), .D(Shift_reg_68_26_1580_i_i_1), 
        .Y(N_65));
    CFG3 #( .INIT(8'h01) )  \State1_ns_0_o5_2_RNI0BC83[0]  (.A(N_2843), 
        .B(\State1_ns_0_o5_2[0]_net_1 ), .C(
        un1_Syn_reg_2_0_a3_RNINA0E1_net_1), .Y(Shift_N_7_1));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[47]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4655), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4652_i_0));
    CFG3 #( .INIT(8'h10) )  Shift_reg_68_13_1953_i_i_N_4L5_N_3L4 (.A(
        N_53_i), .B(\Shift_reg[28]_net_1 ), .C(N_94_i), .Y(
        Shift_reg_68_13_1953_i_i_N_4L5_N_3L4_net_1));
    CFG3 #( .INIT(8'hA8) )  Start_Buff_0_sqmuxa_1 (.A(CCA_NIRQ_c), .B(
        \State1[0]_net_1 ), .C(un1_Start_Buff_1_net_1), .Y(
        Start_Buff_0_sqmuxa_1_net_1));
    CFG2 #( .INIT(4'h4) )  Shift_reg_68_sn_m57_i_o3_RNISOJH_0 (.A(
        \un1_Syn_reg[0] ), .B(\un1_Syn_reg[5] ), .Y(
        \Shift_reg_68_54_e_0[7] ));
    CFG2 #( .INIT(4'hE) )  Parity_16_1089_i_o4_0 (.A(
        \Parity_Counter[1]_net_1 ), .B(\Parity_Counter[2]_net_1 ), .Y(
        N_3721));
    CFG4 #( .INIT(16'hFB40) )  Shift_reg_68_61_754_i_m4_bm (.A(N_102), 
        .B(Shift_reg_68_28_50_4), .C(RX_GPIO0_c), .D(
        \Shift_reg[10]_net_1 ), .Y(Shift_reg_68_61_754_i_m4_bm_net_1));
    CFG4 #( .INIT(16'h0B00) )  \Shift_reg_RNO[23]  (.A(N_1437_mux), .B(
        N_349_1), .C(N_3846), .D(N_3841_i_1), .Y(N_3841_i_0));
    CFG2 #( .INIT(4'h1) )  un1_block_counter_RNIN85F (.A(
        un1_block_counter_net_1), .B(CCA_NIRQ_c), .Y(un1_CCA_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \Bit_Counter_cry[1]  (.A(VCC_net_1), 
        .B(\Bit_Counter[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        Bit_Counter_s_369_FCO), .S(\Bit_Counter_s[1] ), .Y(), .FCO(
        \Bit_Counter_cry[1]_net_1 ));
    CFG4 #( .INIT(16'h0010) )  \State1_ns_0_o5_2_RNIUCKI3[0]  (.A(
        N_2843), .B(\State1_ns_0_o5_2[0]_net_1 ), .C(
        un1_Syn_reg_2_0_a3_RNI6MOJ1_net_1), .D(
        un1_TC_Packet_Counter17_3_net_1), .Y(Shift_N_7_mux_2));
    SLE \TC_Packet_Counter[18]  (.D(\TC_Packet_Counter_s[18] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[18]));
    CFG4 #( .INIT(16'h78F0) )  Shift_reg_68_16_1869_i_m4_am (.A(
        \Shift_reg_68_54_e_0[17] ), .B(Shift_reg_68_54_net_1), .C(
        \Shift_reg[31]_net_1 ), .D(N_53_i), .Y(
        Shift_reg_68_16_1869_i_m4_am_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIRQB93[5]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[5]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Packet_Counter_cry[4] ), .S(
        \TC_Packet_Counter_s[5] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[5] ));
    CFG4 #( .INIT(16'h0002) )  \Shift_reg_RNI2LBF[52]  (.A(
        \Shift_reg[50]_net_1 ), .B(\Shift_reg[41]_net_1 ), .C(
        \Shift_reg[52]_net_1 ), .D(\Shift_reg[1]_net_1 ), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_41));
    CFG4 #( .INIT(16'h4000) )  Shift_reg_68_23_1667_i_i_a2 (.A(N_74), 
        .B(Shift_reg_68_sn_N_84_mux), .C(\Shift_reg[38]_net_1 ), .D(
        N_216), .Y(N_171));
    CFG4 #( .INIT(16'hF737) )  Shift_reg_68_41_1171_i_1 (.A(
        \Shift_reg_5[25]_net_1 ), .B(CCA_NIRQ_c), .C(N_3793), .D(
        Shift_reg_68_41_1171_i_a7_0), .Y(
        Shift_reg_68_41_1171_i_1_net_1));
    CFG3 #( .INIT(8'h35) )  \Bit_Counter_lm_0[0]  (.A(
        \un1_block_counter_4[0]_net_1 ), .B(un14lto0), .C(
        Bit_Counter_3_sqmuxa), .Y(\Bit_Counter_lm[0] ));
    CFG4 #( .INIT(16'hFD20) )  \Shift_reg_68_28[22]  (.A(
        Shift_reg_68_28_34_0_net_1), .B(N_86), .C(RX_GPIO0_c), .D(
        \Shift_reg[22]_net_1 ), .Y(N_92_0));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_25_1609_i_m4_ns (.A(
        Shift_reg_68_25_1609_i_m4_am_net_1), .B(
        Shift_reg_68_25_1609_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4154));
    SLE Flag_once (.D(N_2969_i_0), .CLK(RX_GPIO1_c), .EN(N_88), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Flag_once_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNI156J8[29]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[29]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[28] ), .S(
        \TC_Packet_Counter_s[29] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[29] ));
    CFG4 #( .INIT(16'hF0F4) )  
        Shift_reg_68_0_2328_i_a7_0_0_a3_0_a3_0_a2_1 (.A(
        un1_TC_Packet_Counter17_3_net_1), .B(
        Shift_reg_68_0_2328_i_a7_0_0_a3_0_a3_0_a2_1_1_net_1), .C(
        Shift_reg_68_1_2300_i_0_o2), .D(\State1_ns_0_o5_2[0]_net_1 ), 
        .Y(N_74));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNO[31]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[31]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[30] ), .S(
        \TC_Packet_Counter_s[31] ), .Y(), .FCO());
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[16]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4010), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4007_i_0));
    SLE \Shift_reg[10]  (.D(N_3433_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[10]_net_1 ));
    CFG4 #( .INIT(16'h5551) )  Shift_reg_68_57_866_i_i_0_RNO_1 (.A(
        Shift_reg_68_1_2300_i_0_o2), .B(\State1[0]_net_1 ), .C(
        un1_TC_Packet_Counter17_3_net_1), .D(
        \State1_ns_0_o5_2[0]_net_1 ), .Y(Shift_m8_i_a3_0_sx_0));
    SLE \Shift_reg[37]  (.D(N_4223_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[37]_net_1 ));
    CFG4 #( .INIT(16'hC0EA) )  Shift_reg_68_13_1953_i_i_0 (.A(
        Shift_reg_68_13_1953_i_i_1_tz_net_1), .B(\Shift_reg[28]_net_1 )
        , .C(Shift_reg_68_13_1953_i_i_o3_0_0_net_1), .D(N_74), .Y(
        Shift_reg_68_13_1953_i_i_0_net_1));
    CFG4 #( .INIT(16'hFD20) )  Parity_16_4_431_i_0_m2 (.A(
        \Parity_Counter[0]_net_1 ), .B(Parity_16_5_407_i_o4_0_net_1), 
        .C(RX_GPIO0_c), .D(\Parity[3]_net_1 ), .Y(N_78));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[6]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[6]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[5]_net_1 ), .S(
        \TC_Error_Counter_s[6] ), .Y(), .FCO(
        \TC_Error_Counter_cry[6]_net_1 ));
    CFG2 #( .INIT(4'h7) )  un1_State1_1_0 (.A(
        un1_TC_Packet_Counter17_1_net_1), .B(\State1[0]_net_1 ), .Y(
        un1_State1_1_0_net_1));
    CFG2 #( .INIT(4'h1) )  \State1_ns_0_a5_2_1_0[0]  (.A(
        \Start_Buff[5]_net_1 ), .B(\Start_Buff[6]_net_1 ), .Y(
        un1_Start_Buff_1_5_net_1));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_16_1869_i_m4_ns (.A(
        Shift_reg_68_16_1869_i_m4_am_net_1), .B(
        Shift_reg_68_16_1869_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4367));
    CFG4 #( .INIT(16'h8000) )  \Shift_reg_RNIUFBQ[20]  (.A(
        un1_DataI_0_a3_a_a_a_a_a_a_0_46), .B(
        un1_DataI_0_a3_a_a_a_a_a_a_0_45), .C(
        un1_DataI_0_a3_a_a_a_a_a_a_0_44), .D(
        un1_DataI_0_a3_a_a_a_a_a_a_0_43), .Y(
        un1_DataI_0_a3_a_a_a_a_a_a_0_58));
    CFG3 #( .INIT(8'hAC) )  Shift_reg_68_12_1982_i_m4_ns (.A(
        Shift_reg_68_12_1982_i_m4_bm_net_1), .B(
        Shift_reg_68_12_1982_i_m4_am_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4467));
    CFG3 #( .INIT(8'h20) )  Bit_Counter_3_sqmuxa_0_a2 (.A(N_3002), .B(
        N_277), .C(TC_Packet_Counter17_i_0), .Y(Bit_Counter_3_sqmuxa));
    CFG4 #( .INIT(16'hA900) )  Shift_reg_68_6_2159_i_i_a2_0 (.A(
        \Shift_reg[49]_net_1 ), .B(N_53_i), .C(N_101), .D(N_250), .Y(
        N_232));
    ARI1 #( .INIT(20'h4AA00) )  \Bit_Counter_cry[2]  (.A(VCC_net_1), 
        .B(\Bit_Counter[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \Bit_Counter_cry[1]_net_1 ), .S(\Bit_Counter_s[2] ), .Y(), 
        .FCO(\Bit_Counter_cry[2]_net_1 ));
    SLE \TC_Packet_Counter[4]  (.D(\TC_Packet_Counter_s[4] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[4]));
    ARI1 #( .INIT(20'h48800) )  \Shift_Bit_Counter_cry[1]  (.A(
        VCC_net_1), .B(\un22_DataO_i[1] ), .C(
        \Shift_Bit_Counter_cry_cy_Y[0] ), .D(GND_net_1), .FCI(
        \Shift_Bit_Counter_cry[0]_net_1 ), .S(\Shift_Bit_Counter_s[1] )
        , .Y(), .FCO(\Shift_Bit_Counter_cry[1]_net_1 ));
    CFG2 #( .INIT(4'h7) )  Shift_reg_68_60_782_i_i_o2_2_0 (.A(
        Shift_reg_68_sn_N_16), .B(N_94_i), .Y(
        Shift_reg_68_60_782_i_i_o2_2_0_net_1));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_28_53_0 (.A(
        \Bit_Counter[2]_net_1 ), .B(un14lto0), .C(N_34), .Y(
        Shift_reg_68_28_53_0_net_1));
    SLE \State2[0]  (.D(\State2_9[0] ), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_12_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \State2[0]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_2_2272_i_m4_ns (.A(
        Shift_reg_68_2_2272_i_m4_am_net_1), .B(
        Shift_reg_68_2_2272_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_4705));
    CFG4 #( .INIT(16'hB391) )  DataO_6_53_am (.A(\un22_DataO_i[1] ), 
        .B(DataO_6_53_am_1_1_net_1), .C(\Shift_reg[29]_net_1 ), .D(
        \Shift_reg[25]_net_1 ), .Y(DataO_6_53_am_net_1));
    CFG4 #( .INIT(16'h3337) )  Shift_reg_68_53_953_i_0 (.A(
        \Shift_reg[3]_net_1 ), .B(CCA_NIRQ_c), .C(Shift_reg_68_sn_N_56)
        , .D(N_82), .Y(Shift_reg_68_53_953_i_0_net_1));
    CFG4 #( .INIT(16'h2A3F) )  Shift_reg_68_13_1953_i_i_N_4L5 (.A(
        Shift_N_5), .B(N_253), .C(
        Shift_reg_68_13_1953_i_i_N_4L5_N_4L6_net_1), .D(
        Shift_reg_68_13_1953_i_i_N_4L5_N_5L8_net_1), .Y(
        Shift_reg_68_13_1953_i_i_1));
    CFG4 #( .INIT(16'hAA2A) )  Shift_reg_68_63_697_i_i_a2_0_0 (.A(
        \Shift_reg[12]_net_1 ), .B(Shift_reg_68_sn_N_9), .C(
        \un1_Syn_reg[5] ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_63_697_i_i_a2_0_0_net_1));
    CFG4 #( .INIT(16'h00EC) )  Shift_reg_68_21_1723_i_i_3_0 (.A(
        Shift_reg_68_21_1723_i_i_a2_2_0_net_1), .B(
        Shift_reg_68_21_1723_i_i_a2_1), .C(Shift_reg_68_sn_N_84_mux), 
        .D(N_74), .Y(Shift_reg_68_21_1723_i_i_3_1));
    CFG4 #( .INIT(16'h8000) )  un1_DataO41_22_0_a3_0_4 (.A(
        \un1_Syn_reg[3]_net_1 ), .B(N_370), .C(N_3002), .D(
        un1_DataO41_22_0_a3_0_2), .Y(un1_DataO41_22_0_a3_0_3_net_1));
    SLE \TC_Packet_Counter[29]  (.D(\TC_Packet_Counter_s[29] ), .CLK(
        RX_GPIO1_c), .EN(N_295), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Packet_Counter[29]));
    SLE \Shift_Bit_Counter[4]  (.D(\Shift_Bit_Counter_s[4] ), .CLK(
        RX_GPIO1_c), .EN(Shift_Bit_Countere), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_Bit_Counter[4]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[13]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[13]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[12]_net_1 ), .S(
        \TC_Error_Counter_s[13] ), .Y(), .FCO(
        \TC_Error_Counter_cry[13]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \State1_ns_0_a5_2_4[0]  (.A(
        \Start_Buff[15]_net_1 ), .B(\Start_Buff[14]_net_1 ), .C(
        \Start_Buff[13]_net_1 ), .D(\Start_Buff[11]_net_1 ), .Y(
        \State1_ns_0_a5_2_4[0]_net_1 ));
    CFG2 #( .INIT(4'hD) )  Shift_reg_68_9_2070_i_0_o2_0 (.A(N_53_i), 
        .B(N_109), .Y(N_268));
    CFG4 #( .INIT(16'h1131) )  Shift_reg_68_53_953_i_a7 (.A(
        \State1[0]_net_1 ), .B(\Shift_reg[3]_net_1 ), .C(
        Shift_reg_68_sn_N_73), .D(un1_TC_Packet_Counter17_3_net_1), .Y(
        N_3606));
    CFG3 #( .INIT(8'hCA) )  Shift_reg_68_33_1407_i_m4_ns (.A(
        Shift_reg_68_33_1407_i_m4_am_net_1), .B(
        Shift_reg_68_33_1407_i_m4_bm_net_1), .C(
        Shift_reg_68_sn_N_84_mux), .Y(N_3985));
    CFG4 #( .INIT(16'hF0B8) )  Shift_reg_68_5_2187_i_m4 (.A(N_4629), 
        .B(Shift_reg_68_sn_N_84_mux), .C(\Shift_reg[48]_net_1 ), .D(
        Shift_reg_68_sn_N_56), .Y(N_4630));
    CFG2 #( .INIT(4'h8) )  \Bit_Counter_lm_0[4]  (.A(
        Bit_Counter_3_sqmuxa), .B(\Bit_Counter_s[4] ), .Y(
        \Bit_Counter_lm[4] ));
    CFG3 #( .INIT(8'hFE) )  Shift_reg_68_28_32_a3_0_o3 (.A(un14lto4), 
        .B(\Bit_Counter[2]_net_1 ), .C(\Bit_Counter[3]_net_1 ), .Y(
        N_387));
    CFG4 #( .INIT(16'h0051) )  \Shift_reg_RNO[44]  (.A(N_4727_i_1), .B(
        N_403), .C(\Shift_reg[44]_net_1 ), .D(
        Shift_reg_68_1_2300_i_0_0_net_1), .Y(N_4727_i_0));
    CFG4 #( .INIT(16'h0400) )  Shift_reg_68_7_2129_i_a7_3 (.A(
        Shift_reg_68_sn_N_56), .B(Shift_reg_68_sn_N_84_mux), .C(N_120), 
        .D(N_82), .Y(N_4585));
    CFG4 #( .INIT(16'hF078) )  Shift_reg_68_58_838_i_m4_am (.A(
        \Shift_reg_68_54_e_0[7] ), .B(Shift_reg_68_54_4), .C(
        \Shift_reg[7]_net_1 ), .D(\un1_Syn_reg[6] ), .Y(
        Shift_reg_68_58_838_i_m4_am_net_1));
    CFG3 #( .INIT(8'h5D) )  Block_ErrO_0_sqmuxa_1_0 (.A(
        \State1[0]_net_1 ), .B(TC_Packet_Counter17_i_0), .C(N_277), .Y(
        Block_ErrO_0_sqmuxa_1_0_net_1));
    SLE Block_ErrO (.D(N_74), .CLK(RX_GPIO1_c), .EN(un1_DataO41_27_i_0)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(CLTU_0_Block_ErrO));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Error_Counter_cry[27]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Error_Counter[27]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Error_Counter_cry[26]_net_1 ), .S(
        \TC_Error_Counter_s[27] ), .Y(), .FCO(
        \TC_Error_Counter_cry[27]_net_1 ));
    CFG4 #( .INIT(16'hA280) )  Start_Buff_0_sqmuxa_0_0 (.A(CCA_NIRQ_c), 
        .B(\State1[0]_net_1 ), .C(TC_Packet_Counter17_i_0), .D(
        un1_Start_Buff_1_net_1), .Y(Start_Buff_0_sqmuxa_0_0_net_1));
    CFG3 #( .INIT(8'hC6) )  \Shift_reg_RNO_0[23]  (.A(
        Shift_reg_68_50_5), .B(\Shift_reg[23]_net_1 ), .C(
        \un1_Syn_reg[6] ), .Y(N_1437_mux));
    CFG4 #( .INIT(16'h40C0) )  \Shift_reg_RNO[29]  (.A(
        \State1[0]_net_1 ), .B(CCA_NIRQ_c), .C(N_4417), .D(
        un1_TC_Packet_Counter17_5_net_1), .Y(N_4414_i_0));
    SLE \TC_Error_Counter[31]  (.D(\TC_Error_Counter_s[31]_net_1 ), 
        .CLK(RX_GPIO1_c), .EN(N_79_i_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CLTU_0_TC_Error_Counter[31]));
    CFG4 #( .INIT(16'h0080) )  Shift_reg_68_28_24_0 (.A(un14lto0), .B(
        \State1[0]_net_1 ), .C(N_290), .D(N_58), .Y(
        Shift_reg_68_28_50_4));
    CFG4 #( .INIT(16'h0004) )  Shift_reg_68_28_2 (.A(N_265), .B(
        \Bit_Counter[3]_net_1 ), .C(N_57), .D(N_385), .Y(
        Shift_reg_68_28_2_net_1));
    CFG3 #( .INIT(8'h9A) )  Shift_reg_68_3_2244_i_m4_am (.A(
        \Shift_reg[46]_net_1 ), .B(\un1_Syn_reg[5] ), .C(N_1461), .Y(
        Shift_reg_68_3_2244_i_m4_am_net_1));
    CFG3 #( .INIT(8'h9A) )  Shift_reg_68_18_1811_i_m4_am (.A(
        \Shift_reg[33]_net_1 ), .B(\un1_Syn_reg[0] ), .C(N_1445), .Y(
        Shift_reg_68_18_1811_i_m4_am_net_1));
    SLE \Shift_reg[31]  (.D(N_4364_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[31]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \State1_ns_0_a5_2_6_0[0]  (.A(
        \Start_Buff[8]_net_1 ), .B(\Start_Buff[7]_net_1 ), .C(N_2131_1)
        , .Y(\State1_ns_0_a5_2_6[0] ));
    SLE \Shift_reg[40]  (.D(N_4151_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[40]_net_1 ));
    CFG4 #( .INIT(16'h3F15) )  \Shift_reg_RNO_0[19]  (.A(N_349_1), .B(
        un1_TC_Packet_Counter17_5_net_1), .C(\State1[0]_net_1 ), .D(
        N_1450_mux), .Y(N_3935_i_1));
    CFG4 #( .INIT(16'h3337) )  Shift_reg_68_20_1753_i_0 (.A(
        \Shift_reg[35]_net_1 ), .B(CCA_NIRQ_c), .C(
        Shift_reg_68_sn_N_56), .D(N_82), .Y(
        Shift_reg_68_20_1753_i_0_net_1));
    CFG2 #( .INIT(4'h2) )  un1_DataO41_24_i_a3_0_1 (.A(un14lto5), .B(
        Flag_once_net_1), .Y(N_356_1));
    CFG4 #( .INIT(16'hB4F0) )  \Shift_reg_RNO_1[19]  (.A(
        \un1_Syn_reg[0] ), .B(Shift_reg_68_50_net_1), .C(
        \Shift_reg[19]_net_1 ), .D(\un1_Syn_reg[5] ), .Y(N_1450_mux));
    SLE \Parity[5]  (.D(N_3720_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_10_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Parity[5]_net_1 ));
    CFG4 #( .INIT(16'h159D) )  DataO_10_iv_0_0_RNO_23 (.A(
        \un22_DataO_i[2] ), .B(\Shift_Bit_Counter[5]_net_1 ), .C(
        \Shift_reg[20]_net_1 ), .D(\Shift_reg[16]_net_1 ), .Y(
        DataO_6_13_i_m2_1_2));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_8_2099_i_0_a3_2 (.A(
        Shift_reg_68_sn_N_56), .B(\Shift_reg[51]_net_1 ), .C(N_82), .Y(
        N_350));
    CFG4 #( .INIT(16'hAAA6) )  \Shift_reg_68_44[48]  (.A(
        \Shift_reg[48]_net_1 ), .B(Shift_reg_68_sn_N_9), .C(
        \un1_Syn_reg[5] ), .D(\un1_Syn_reg[6] ), .Y(N_206));
    CFG3 #( .INIT(8'h01) )  Shift_reg_68_31_1463_i_a7_2 (.A(
        Shift_reg_68_sn_N_56), .B(\Shift_reg[15]_net_1 ), .C(N_82), .Y(
        N_4036));
    CFG4 #( .INIT(16'h8F83) )  DataO_10_iv_0_0_RNO_0 (.A(N_314), .B(
        \un22_DataO_i[0] ), .C(DataO_6_46_1_2), .D(N_2673), .Y(N_2675));
    CFG2 #( .INIT(4'h1) )  Shift_reg_68_28_34_0 (.A(N_387), .B(N_102), 
        .Y(Shift_reg_68_28_34_0_net_1));
    SLE \Shift_reg[54]  (.D(N_4489_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_DataO41_22_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Shift_reg[54]_net_1 ));
    CFG4 #( .INIT(16'h0FEF) )  un1_DataI_0_a3_a_a_a_a_a_a_RNI1ARV (.A(
        \State1_ns_0_o5_2[0]_net_1 ), .B(\State1_ns_0_o5_3[0]_net_1 ), 
        .C(\State1[0]_net_1 ), .D(un1_DataI), .Y(un1_DataO41_26_i_1));
    CFG4 #( .INIT(16'h8F83) )  DataO_10_iv_0_0_RNO_5 (.A(N_400), .B(
        \un22_DataO_i[0] ), .C(DataO_6_30_1_2), .D(N_340), .Y(N_2659));
    CFG3 #( .INIT(8'h06) )  \block_counter_8[0]  (.A(
        \block_counter[0]_net_1 ), .B(\un1_block_counter_4[0]_net_1 ), 
        .C(\un1_block_counter_7[0] ), .Y(\block_counter_8[0]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNIU8VO8[30]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[30]), .C(GND_net_1), 
        .D(GND_net_1), .FCI(\TC_Packet_Counter_cry[29] ), .S(
        \TC_Packet_Counter_s[30] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[30] ));
    ARI1 #( .INIT(20'h4AA00) )  \TC_Packet_Counter_RNICMJR2[4]  (.A(
        VCC_net_1), .B(CLTU_0_TC_Packet_Counter[4]), .C(GND_net_1), .D(
        GND_net_1), .FCI(\TC_Packet_Counter_cry[3] ), .S(
        \TC_Packet_Counter_s[4] ), .Y(), .FCO(
        \TC_Packet_Counter_cry[4] ));
    CFG3 #( .INIT(8'h04) )  Shift_reg_68_28_14_2 (.A(
        \Bit_Counter[3]_net_1 ), .B(un14lto4), .C(un14lto5), .Y(
        Shift_reg_68_28_14_1));
    
endmodule


module TM_RSENC_TM_RSENC_0_kitCountS_8s_253s_1s(
       Bit_Count_16dec_i_1,
       Q_cry_cy_Y,
       timer_w_0,
       timer_w_1,
       timer_w_5,
       RSControl_0_NGRST,
       RSControl_0_START,
       TM_RSENC_0_RDY,
       N_1419,
       dataOver_w
    );
input  [3:3] Bit_Count_16dec_i_1;
output [0:0] Q_cry_cy_Y;
output timer_w_0;
output timer_w_1;
output timer_w_5;
input  RSControl_0_NGRST;
input  RSControl_0_START;
input  TM_RSENC_0_RDY;
output N_1419;
output dataOver_w;

    wire VCC_net_1, \Q_s[0] , GND_net_1, \Q_s[1] , \timer_w[2] , 
        \Q_s[2] , \timer_w[3] , \Q_s[3] , \timer_w[4] , \Q_s[4] , 
        \Q_s[5] , \timer_w[6] , \Q_s[6] , \timer_w[7] , \Q_s[7]_net_1 , 
        Q_cry_cy, \Q_cry[0]_net_1 , \Q_cry[1]_net_1 , \Q_cry[2]_net_1 , 
        \Q_cry[3]_net_1 , \Q_cry[4]_net_1 , \Q_cry[5]_net_1 , 
        \Q_cry[6]_net_1 , G_6_0_a2_1, G_6_0_a2_0_1;
    
    SLE \Q[6]  (.D(\Q_s[6] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\timer_w[6] ));
    CFG2 #( .INIT(4'h2) )  \Q_RNILV8J[5]  (.A(TM_RSENC_0_RDY), .B(
        timer_w_5), .Y(G_6_0_a2_1));
    CFG4 #( .INIT(16'h8000) )  \Q_RNIMV071[3]  (.A(\timer_w[7] ), .B(
        \timer_w[4] ), .C(\timer_w[3] ), .D(G_6_0_a2_0_1), .Y(N_1419));
    SLE \Q[2]  (.D(\Q_s[2] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\timer_w[2] ));
    GND GND (.Y(GND_net_1));
    SLE \Q[4]  (.D(\Q_s[4] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\timer_w[4] ));
    ARI1 #( .INIT(20'h44400) )  \Q_cry[2]  (.A(VCC_net_1), .B(
        RSControl_0_START), .C(\timer_w[2] ), .D(GND_net_1), .FCI(
        \Q_cry[1]_net_1 ), .S(\Q_s[2] ), .Y(), .FCO(\Q_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h44400) )  \Q_cry[0]  (.A(VCC_net_1), .B(
        RSControl_0_START), .C(timer_w_0), .D(GND_net_1), .FCI(
        Q_cry_cy), .S(\Q_s[0] ), .Y(), .FCO(\Q_cry[0]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  \Q_RNICAT92[0]  (.A(timer_w_1), .B(
        timer_w_0), .C(N_1419), .D(G_6_0_a2_1), .Y(dataOver_w));
    ARI1 #( .INIT(20'h44400) )  \Q_s[7]  (.A(VCC_net_1), .B(
        RSControl_0_START), .C(\timer_w[7] ), .D(GND_net_1), .FCI(
        \Q_cry[6]_net_1 ), .S(\Q_s[7]_net_1 ), .Y(), .FCO());
    ARI1 #( .INIT(20'h44400) )  \Q_cry[3]  (.A(VCC_net_1), .B(
        RSControl_0_START), .C(\timer_w[3] ), .D(GND_net_1), .FCI(
        \Q_cry[2]_net_1 ), .S(\Q_s[3] ), .Y(), .FCO(\Q_cry[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \Q_RNI8IJF[2]  (.A(\timer_w[2] ), .B(
        \timer_w[6] ), .Y(G_6_0_a2_0_1));
    ARI1 #( .INIT(20'h44400) )  \Q_cry[6]  (.A(VCC_net_1), .B(
        RSControl_0_START), .C(\timer_w[6] ), .D(GND_net_1), .FCI(
        \Q_cry[5]_net_1 ), .S(\Q_s[6] ), .Y(), .FCO(\Q_cry[6]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  \Q_cry_cy[0]  (.A(VCC_net_1), .B(
        RSControl_0_START), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(Q_cry_cy_Y[0]), .FCO(Q_cry_cy));
    SLE \Q[3]  (.D(\Q_s[3] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\timer_w[3] ));
    SLE \Q[7]  (.D(\Q_s[7]_net_1 ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\timer_w[7] ));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h44400) )  \Q_cry[4]  (.A(VCC_net_1), .B(
        RSControl_0_START), .C(\timer_w[4] ), .D(GND_net_1), .FCI(
        \Q_cry[3]_net_1 ), .S(\Q_s[4] ), .Y(), .FCO(\Q_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h44400) )  \Q_cry[1]  (.A(VCC_net_1), .B(
        RSControl_0_START), .C(timer_w_1), .D(GND_net_1), .FCI(
        \Q_cry[0]_net_1 ), .S(\Q_s[1] ), .Y(), .FCO(\Q_cry[1]_net_1 ));
    SLE \Q[1]  (.D(\Q_s[1] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(timer_w_1));
    SLE \Q[0]  (.D(\Q_s[0] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(timer_w_0));
    SLE \Q[5]  (.D(\Q_s[5] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(timer_w_5));
    ARI1 #( .INIT(20'h44400) )  \Q_cry[5]  (.A(VCC_net_1), .B(
        RSControl_0_START), .C(timer_w_5), .D(GND_net_1), .FCI(
        \Q_cry[4]_net_1 ), .S(\Q_s[5] ), .Y(), .FCO(\Q_cry[5]_net_1 ));
    
endmodule


module TM_RSENC_TM_RSENC_0_kitDelay_bit_reg_4s(
       Bit_Count_16dec_i_1,
       TM_RSENC_0_RDY,
       RSControl_0_NGRST,
       pre_rdy
    );
input  [3:3] Bit_Count_16dec_i_1;
output TM_RSENC_0_RDY;
input  RSControl_0_NGRST;
input  pre_rdy;

    wire VCC_net_1, \delayLine_2_[0] , GND_net_1, \delayLine_1_[0] , 
        \delayLine_0_[0] ;
    
    SLE \genblk1.delayLine_0_[0]  (.D(pre_rdy), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\delayLine_0_[0] ));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    SLE \genblk1.delayLine_1_[0]  (.D(\delayLine_0_[0] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\delayLine_1_[0] ));
    SLE \genblk1.delayLine_3_[0]  (.D(\delayLine_2_[0] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(TM_RSENC_0_RDY));
    SLE \genblk1.delayLine_2_[0]  (.D(\delayLine_1_[0] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\delayLine_2_[0] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_SM_223s_16s_255s_8s_1s_1s_4s(
       Bit_Count_16dec_i_1,
       hold0fb_w,
       TM_RSENC_0_RFD,
       RSControl_0_NGRST,
       TM_RSENC_0_RFS,
       datNotParity_w,
       RSControl_0_START,
       TM_RSENC_0_RDY
    );
input  [3:3] Bit_Count_16dec_i_1;
output hold0fb_w;
output TM_RSENC_0_RFD;
input  RSControl_0_NGRST;
output TM_RSENC_0_RFS;
output datNotParity_w;
input  RSControl_0_START;
output TM_RSENC_0_RDY;

    wire hold0fb_w_i_0, GND_net_1, rfd_2_sqmuxa_i_0_net_1, VCC_net_1, 
        hold0fb_r_net_1, dataOver_w, hold0fb_r_2_sqmuxa_i_0_net_1, 
        pre_rdy_net_1, N_1285_i_0, un1_valid_start_1_net_1, 
        \Q_cry_cy_Y[0] , un1_start_2_0_net_1, codeOver_net_1, 
        codeOver_2, \timer_w[0] , \timer_w[5] , N_1348_1, \timer_w[1] , 
        N_1419;
    
    SLE hold0fb_r (.D(dataOver_w), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        hold0fb_r_2_sqmuxa_i_0_net_1), .ALn(RSControl_0_NGRST), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(hold0fb_r_net_1));
    GND GND (.Y(GND_net_1));
    SLE codeOver (.D(codeOver_2), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(codeOver_net_1)
        );
    CFG3 #( .INIT(8'hF8) )  un1_valid_start_1 (.A(RSControl_0_START), 
        .B(TM_RSENC_0_RFS), .C(codeOver_net_1), .Y(
        un1_valid_start_1_net_1));
    SLE pre_rdy (.D(N_1285_i_0), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        un1_valid_start_1_net_1), .ALn(RSControl_0_NGRST), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(pre_rdy_net_1));
    CFG1 #( .INIT(2'h1) )  datNotParity_RNO (.A(hold0fb_w), .Y(
        hold0fb_w_i_0));
    TM_RSENC_TM_RSENC_0_kitCountS_8s_253s_1s sm_timer_0 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .Q_cry_cy_Y({
        \Q_cry_cy_Y[0] }), .timer_w_0(\timer_w[0] ), .timer_w_1(
        \timer_w[1] ), .timer_w_5(\timer_w[5] ), .RSControl_0_NGRST(
        RSControl_0_NGRST), .RSControl_0_START(RSControl_0_START), 
        .TM_RSENC_0_RDY(TM_RSENC_0_RDY), .N_1419(N_1419), .dataOver_w(
        dataOver_w));
    SLE rfs (.D(\Q_cry_cy_Y[0] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        un1_start_2_0_net_1), .ALn(RSControl_0_NGRST), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TM_RSENC_0_RFS));
    SLE rfd (.D(TM_RSENC_0_RFS), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        rfd_2_sqmuxa_i_0_net_1), .ALn(RSControl_0_NGRST), .ADn(
        GND_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(TM_RSENC_0_RFD));
    CFG2 #( .INIT(4'h8) )  codeOver_2_0_a2_1 (.A(\timer_w[0] ), .B(
        \timer_w[5] ), .Y(N_1348_1));
    CFG4 #( .INIT(16'h4000) )  codeOver_2_0_a2 (.A(\timer_w[1] ), .B(
        N_1348_1), .C(TM_RSENC_0_RDY), .D(N_1419), .Y(codeOver_2));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'hE) )  rfd_2_sqmuxa_i_0 (.A(dataOver_w), .B(
        TM_RSENC_0_RFS), .Y(rfd_2_sqmuxa_i_0_net_1));
    CFG2 #( .INIT(4'h8) )  pre_rdy_RNO (.A(TM_RSENC_0_RFS), .B(
        RSControl_0_START), .Y(N_1285_i_0));
    CFG4 #( .INIT(16'hBAAA) )  un1_start_2_0 (.A(RSControl_0_START), 
        .B(\timer_w[1] ), .C(N_1419), .D(N_1348_1), .Y(
        un1_start_2_0_net_1));
    TM_RSENC_TM_RSENC_0_kitDelay_bit_reg_4s bit_dly_0 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), 
        .TM_RSENC_0_RDY(TM_RSENC_0_RDY), .RSControl_0_NGRST(
        RSControl_0_NGRST), .pre_rdy(pre_rdy_net_1));
    CFG2 #( .INIT(4'hE) )  hold0fb_r_2_sqmuxa_i_0 (.A(dataOver_w), .B(
        RSControl_0_START), .Y(hold0fb_r_2_sqmuxa_i_0_net_1));
    SLE hold0fb_r2 (.D(hold0fb_r_net_1), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(hold0fb_w));
    SLE datNotParity (.D(hold0fb_w_i_0), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(datNotParity_w)
        );
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_165s_8s(
       Bit_Count_16dec_i_1,
       shft9_w,
       shft8_w,
       fb_w_1,
       fb_w_5,
       fb_w_7,
       fb_w_2,
       fb_w_0,
       fb_w_4,
       fb_w_3,
       RSControl_0_NGRST,
       N_566,
       N_568,
       N_574,
       N_564,
       N_570,
       N_567,
       N_565,
       N_588
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft9_w;
input  [7:0] shft8_w;
input  fb_w_1;
input  fb_w_5;
input  fb_w_7;
input  fb_w_2;
input  fb_w_0;
input  fb_w_4;
input  fb_w_3;
input  RSControl_0_NGRST;
input  N_566;
input  N_568;
input  N_574;
input  N_564;
input  N_570;
input  N_567;
input  N_565;
input  N_588;

    wire VCC_net_1, \shftOut_29[3] , GND_net_1, \shftOut_29[4] , 
        \shftOut_29[5] , \shftOut_29[6] , \shftOut_29[7] , 
        \shftOut_29[0] , \shftOut_29[1] , \shftOut_29[2] ;
    
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[5]  (.A(shft8_w[5]), 
        .B(fb_w_4), .C(N_588), .D(N_565), .Y(\shftOut_29[5] ));
    SLE \shftOut[5]  (.D(\shftOut_29[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft9_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_29[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft9_w[6]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[3]  (.A(fb_w_2), .B(
        shft8_w[3]), .C(N_567), .D(N_565), .Y(\shftOut_29[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_29_0_a2[0]  (.A(shft8_w[0]), .B(
        N_574), .C(N_564), .Y(\shftOut_29[0] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_29[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft9_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_29_0_a2[1]  (.A(shft8_w[1]), .B(
        fb_w_7), .C(N_568), .Y(\shftOut_29[1] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[4]  (.A(shft8_w[4]), 
        .B(fb_w_2), .C(fb_w_3), .D(N_566), .Y(\shftOut_29[4] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[6]  (.A(shft8_w[6]), 
        .B(fb_w_1), .C(fb_w_5), .D(N_566), .Y(\shftOut_29[6] ));
    SLE \shftOut[7]  (.D(\shftOut_29[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft9_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_29[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft9_w[3]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[2]  (.A(shft8_w[2]), 
        .B(fb_w_7), .C(fb_w_1), .D(N_570), .Y(\shftOut_29[2] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[7]  (.A(shft8_w[7]), 
        .B(fb_w_0), .C(fb_w_1), .D(N_565), .Y(\shftOut_29[7] ));
    SLE \shftOut[2]  (.D(\shftOut_29[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft9_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_29[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft9_w[1]));
    SLE \shftOut[0]  (.D(\shftOut_29[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft9_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_86s_8s_2(
       Bit_Count_16dec_i_1,
       shft29_w,
       shft28_w,
       fb_w,
       RSControl_0_NGRST,
       N_568,
       N_567,
       N_574,
       N_569,
       N_576,
       N_564,
       N_565,
       N_570,
       N_575
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft29_w;
input  [7:0] shft28_w;
input  [7:1] fb_w;
input  RSControl_0_NGRST;
input  N_568;
input  N_567;
input  N_574;
input  N_569;
input  N_576;
input  N_564;
input  N_565;
input  N_570;
input  N_575;

    wire VCC_net_1, \shftOut_11[3] , GND_net_1, \shftOut_11[4] , 
        \shftOut_11[5] , \shftOut_11[6] , \shftOut_11[7] , 
        \shftOut_11[0] , \shftOut_11[1] , \shftOut_11[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_11[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft29_w[5]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[3]  (.A(shft28_w[3]), 
        .B(fb_w[2]), .C(fb_w[6]), .D(N_575), .Y(\shftOut_11[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[2]  (.A(shft28_w[2]), .B(
        N_574), .C(N_569), .Y(\shftOut_11[2] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[6]  (.A(shft28_w[6]), .B(
        fb_w[5]), .C(N_570), .Y(\shftOut_11[6] ));
    SLE \shftOut[6]  (.D(\shftOut_11[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft29_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_11[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft29_w[4]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[7]  (.A(shft28_w[7]), 
        .B(fb_w[2]), .C(fb_w[1]), .D(N_565), .Y(\shftOut_11[7] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[5]  (.A(shft28_w[5]), 
        .B(fb_w[4]), .C(fb_w[5]), .D(N_567), .Y(\shftOut_11[5] ));
    SLE \shftOut[7]  (.D(\shftOut_11[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft29_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_11[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft29_w[3]));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[1]  (.A(shft28_w[1]), .B(
        fb_w[7]), .C(N_570), .Y(\shftOut_11[1] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[0]  (.A(shft28_w[0]), .B(
        fb_w[2]), .C(N_568), .Y(\shftOut_11[0] ));
    SLE \shftOut[2]  (.D(\shftOut_11[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft29_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_11[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft29_w[1]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[4]  (.A(shft28_w[4]), 
        .B(fb_w[3]), .C(N_576), .D(N_564), .Y(\shftOut_11[4] ));
    SLE \shftOut[0]  (.D(\shftOut_11[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft29_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_86s_8s_1(
       Bit_Count_16dec_i_1,
       shft19_w,
       shft18_w,
       fb_w,
       RSControl_0_NGRST,
       N_568,
       N_567,
       N_574,
       N_569,
       N_576,
       N_564,
       N_565,
       N_570,
       N_575
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft19_w;
input  [7:0] shft18_w;
input  [7:1] fb_w;
input  RSControl_0_NGRST;
input  N_568;
input  N_567;
input  N_574;
input  N_569;
input  N_576;
input  N_564;
input  N_565;
input  N_570;
input  N_575;

    wire VCC_net_1, \shftOut_11[3] , GND_net_1, \shftOut_11[4] , 
        \shftOut_11[5] , \shftOut_11[6] , \shftOut_11[7] , 
        \shftOut_11[0] , \shftOut_11[1] , \shftOut_11[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_11[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft19_w[5]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[3]  (.A(shft18_w[3]), 
        .B(fb_w[2]), .C(fb_w[6]), .D(N_575), .Y(\shftOut_11[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[2]  (.A(shft18_w[2]), .B(
        N_574), .C(N_569), .Y(\shftOut_11[2] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[6]  (.A(shft18_w[6]), .B(
        fb_w[5]), .C(N_570), .Y(\shftOut_11[6] ));
    SLE \shftOut[6]  (.D(\shftOut_11[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft19_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_11[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft19_w[4]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[7]  (.A(shft18_w[7]), 
        .B(fb_w[2]), .C(fb_w[1]), .D(N_565), .Y(\shftOut_11[7] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[5]  (.A(shft18_w[5]), 
        .B(fb_w[4]), .C(fb_w[5]), .D(N_567), .Y(\shftOut_11[5] ));
    SLE \shftOut[7]  (.D(\shftOut_11[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft19_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_11[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft19_w[3]));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[1]  (.A(shft18_w[1]), .B(
        fb_w[7]), .C(N_570), .Y(\shftOut_11[1] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[0]  (.A(shft18_w[0]), .B(
        fb_w[2]), .C(N_568), .Y(\shftOut_11[0] ));
    SLE \shftOut[2]  (.D(\shftOut_11[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft19_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_11[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft19_w[1]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[4]  (.A(shft18_w[4]), 
        .B(fb_w[3]), .C(N_576), .D(N_564), .Y(\shftOut_11[4] ));
    SLE \shftOut[0]  (.D(\shftOut_11[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft19_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_86s_8s(
       Bit_Count_16dec_i_1,
       shft3_w,
       shft2_w,
       fb_w,
       RSControl_0_NGRST,
       N_568,
       N_567,
       N_574,
       N_569,
       N_576,
       N_564,
       N_565,
       N_570,
       N_575
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft3_w;
input  [7:0] shft2_w;
input  [7:1] fb_w;
input  RSControl_0_NGRST;
input  N_568;
input  N_567;
input  N_574;
input  N_569;
input  N_576;
input  N_564;
input  N_565;
input  N_570;
input  N_575;

    wire VCC_net_1, \shftOut_11[3] , GND_net_1, \shftOut_11[4] , 
        \shftOut_11[5] , \shftOut_11[6] , \shftOut_11[7] , 
        \shftOut_11[0] , \shftOut_11[1] , \shftOut_11[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_11[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft3_w[5]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[3]  (.A(shft2_w[3]), 
        .B(fb_w[2]), .C(fb_w[6]), .D(N_575), .Y(\shftOut_11[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[2]  (.A(shft2_w[2]), .B(
        N_574), .C(N_569), .Y(\shftOut_11[2] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[6]  (.A(shft2_w[6]), .B(
        fb_w[5]), .C(N_570), .Y(\shftOut_11[6] ));
    SLE \shftOut[6]  (.D(\shftOut_11[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft3_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_11[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft3_w[4]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[7]  (.A(shft2_w[7]), 
        .B(fb_w[2]), .C(fb_w[1]), .D(N_565), .Y(\shftOut_11[7] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[5]  (.A(shft2_w[5]), 
        .B(fb_w[4]), .C(fb_w[5]), .D(N_567), .Y(\shftOut_11[5] ));
    SLE \shftOut[7]  (.D(\shftOut_11[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft3_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_11[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft3_w[3]));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[1]  (.A(shft2_w[1]), .B(
        fb_w[7]), .C(N_570), .Y(\shftOut_11[1] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[0]  (.A(shft2_w[0]), .B(
        fb_w[2]), .C(N_568), .Y(\shftOut_11[0] ));
    SLE \shftOut[2]  (.D(\shftOut_11[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft3_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_11[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft3_w[1]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[4]  (.A(shft2_w[4]), 
        .B(fb_w[3]), .C(N_576), .D(N_564), .Y(\shftOut_11[4] ));
    SLE \shftOut[0]  (.D(\shftOut_11[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft3_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_30s_8s_0(
       Bit_Count_16dec_i_1,
       shft27_w,
       pre_fb_w,
       dInp_reg_w,
       shftOut_17_1,
       shft26_w,
       fb_w_0,
       fb_w_7,
       fb_w_1,
       fb_w_5,
       fb_w_3,
       fb_w_4,
       fb_w_6,
       RSControl_0_NGRST,
       N_566,
       N_565,
       N_575,
       N_572,
       N_574,
       N_564
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft27_w;
input  [3:3] pre_fb_w;
input  [3:3] dInp_reg_w;
output [2:2] shftOut_17_1;
input  [7:0] shft26_w;
input  fb_w_0;
input  fb_w_7;
input  fb_w_1;
input  fb_w_5;
input  fb_w_3;
input  fb_w_4;
input  fb_w_6;
input  RSControl_0_NGRST;
input  N_566;
input  N_565;
output N_575;
input  N_572;
input  N_574;
input  N_564;

    wire VCC_net_1, \shftOut_17[3] , GND_net_1, \shftOut_17[4] , 
        \shftOut_17[5] , \shftOut_17[6] , \shftOut_17[7] , 
        \shftOut_17[0] , \shftOut_17[1] , \shftOut_17[2] ;
    
    CFG4 #( .INIT(16'h6996) )  \shftOut_17_0_a2[6]  (.A(shft26_w[6]), 
        .B(fb_w_3), .C(fb_w_5), .D(N_572), .Y(\shftOut_17[6] ));
    SLE \shftOut[5]  (.D(\shftOut_17[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft27_w[5]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_17_0_a2_1[2]  (.A(fb_w_4), .B(
        fb_w_0), .C(fb_w_1), .D(N_565), .Y(shftOut_17_1[2]));
    SLE \shftOut[6]  (.D(\shftOut_17[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft27_w[6]));
    CFG3 #( .INIT(8'h96) )  \shftOut_17_0_a2[7]  (.A(fb_w_5), .B(
        shft26_w[7]), .C(fb_w_3), .Y(\shftOut_17[7] ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h96) )  \shftOut_17_0_a2[5]  (.A(N_575), .B(
        shft26_w[5]), .C(N_572), .Y(\shftOut_17[5] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_17_0_a2_0[5]  (.A(fb_w_7), .B(
        fb_w_1), .C(pre_fb_w[3]), .D(dInp_reg_w[3]), .Y(N_575));
    SLE \shftOut[4]  (.D(\shftOut_17[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft27_w[4]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_17_0_a2[1]  (.A(shft26_w[1]), 
        .B(fb_w_0), .C(N_566), .D(N_565), .Y(\shftOut_17[1] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_17_0_a2[0]  (.A(N_566), .B(
        shft26_w[0]), .Y(\shftOut_17[0] ));
    SLE \shftOut[7]  (.D(\shftOut_17[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft27_w[7]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_17_0_a2[4]  (.A(shft26_w[4]), 
        .B(fb_w_6), .C(N_575), .D(N_564), .Y(\shftOut_17[4] ));
    SLE \shftOut[3]  (.D(\shftOut_17[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft27_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_17[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft27_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_17[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft27_w[1]));
    SLE \shftOut[0]  (.D(\shftOut_17[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft27_w[0]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_17_0_a2[3]  (.A(shft26_w[3]), 
        .B(fb_w_5), .C(N_574), .D(N_564), .Y(\shftOut_17[3] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_17_0_a2[2]  (.A(shftOut_17_1[2]), 
        .B(shft26_w[2]), .Y(\shftOut_17[2] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_32s_8s_0(
       Bit_Count_16dec_i_1,
       shft17_w,
       shft16_w,
       fb_w_3,
       fb_w_6,
       fb_w_0,
       fb_w_7,
       fb_w_1,
       fb_w_2,
       RSControl_0_NGRST,
       N_566,
       N_565,
       N_568,
       N_573
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft17_w;
input  [7:0] shft16_w;
input  fb_w_3;
input  fb_w_6;
input  fb_w_0;
input  fb_w_7;
input  fb_w_1;
input  fb_w_2;
input  RSControl_0_NGRST;
input  N_566;
input  N_565;
input  N_568;
input  N_573;

    wire VCC_net_1, \shftOut_44[3] , GND_net_1, \shftOut_44[4] , 
        \shftOut_44[5] , \shftOut_44[6] , \shftOut_44[7] , 
        \shftOut_44[0] , \shftOut_44[1] , \shftOut_44[2] ;
    
    CFG2 #( .INIT(4'h6) )  \shftOut_44_0_a2[1]  (.A(fb_w_3), .B(
        shft16_w[1]), .Y(\shftOut_44[1] ));
    SLE \shftOut[5]  (.D(\shftOut_44[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft17_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_44[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft17_w[6]));
    CFG3 #( .INIT(8'h96) )  \shftOut_44_0_a2[6]  (.A(shft16_w[6]), .B(
        fb_w_7), .C(fb_w_1), .Y(\shftOut_44[6] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_44[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft17_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_44_0_a2[2]  (.A(shft16_w[2]), .B(
        N_568), .C(N_565), .Y(\shftOut_44[2] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_44_0_a2[3]  (.A(shft16_w[3]), .B(
        fb_w_7), .C(N_566), .Y(\shftOut_44[3] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_44_0_a2[0]  (.A(shft16_w[0]), 
        .B(fb_w_3), .C(N_566), .D(N_565), .Y(\shftOut_44[0] ));
    SLE \shftOut[7]  (.D(\shftOut_44[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft17_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_44[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft17_w[3]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_44_0_a2[7]  (.A(shft16_w[7]), 
        .B(fb_w_2), .C(fb_w_3), .D(N_573), .Y(\shftOut_44[7] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_44_0_a2[4]  (.A(N_565), .B(
        shft16_w[4]), .Y(\shftOut_44[4] ));
    SLE \shftOut[2]  (.D(\shftOut_44[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft17_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_44[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft17_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_44_0_a2[5]  (.A(fb_w_6), .B(
        shft16_w[5]), .C(fb_w_0), .Y(\shftOut_44[5] ));
    SLE \shftOut[0]  (.D(\shftOut_44[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft17_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_16s_8s_0(
       Bit_Count_16dec_i_1,
       shft28_w,
       shft27_w,
       fb_w_3,
       fb_w_4,
       fb_w_2,
       fb_w_6,
       fb_w_0,
       fb_w_7,
       fb_w_1,
       RSControl_0_NGRST,
       N_566,
       N_565,
       N_573
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft28_w;
input  [7:0] shft27_w;
input  fb_w_3;
input  fb_w_4;
input  fb_w_2;
input  fb_w_6;
input  fb_w_0;
input  fb_w_7;
input  fb_w_1;
input  RSControl_0_NGRST;
input  N_566;
input  N_565;
output N_573;

    wire VCC_net_1, \shftOut_14[3] , GND_net_1, \shftOut_14[4] , 
        \shftOut_14[5] , \shftOut_14[6] , \shftOut_14[7] , 
        \shftOut_14[0] , \shftOut_14[1] , \shftOut_14[2] ;
    
    CFG2 #( .INIT(4'h6) )  \shftOut_14_0_a2_0[0]  (.A(N_565), .B(N_566)
        , .Y(N_573));
    SLE \shftOut[5]  (.D(\shftOut_14[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft28_w[5]));
    CFG2 #( .INIT(4'h6) )  \shftOut_14_0_a2[1]  (.A(fb_w_4), .B(
        shft27_w[1]), .Y(\shftOut_14[1] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_14_0_a2[0]  (.A(shft27_w[0]), .B(
        N_566), .C(N_565), .Y(\shftOut_14[0] ));
    SLE \shftOut[6]  (.D(\shftOut_14[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft28_w[6]));
    CFG3 #( .INIT(8'h96) )  \shftOut_14_0_a2[4]  (.A(fb_w_6), .B(
        shft27_w[4]), .C(fb_w_0), .Y(\shftOut_14[4] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_14[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft28_w[4]));
    CFG2 #( .INIT(4'h6) )  \shftOut_14_0_a2[3]  (.A(N_565), .B(
        shft27_w[3]), .Y(\shftOut_14[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_14_0_a2[2]  (.A(shft27_w[2]), .B(
        fb_w_7), .C(N_566), .Y(\shftOut_14[2] ));
    SLE \shftOut[7]  (.D(\shftOut_14[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft28_w[7]));
    CFG2 #( .INIT(4'h6) )  \shftOut_14_0_a2[6]  (.A(fb_w_2), .B(
        shft27_w[6]), .Y(\shftOut_14[6] ));
    SLE \shftOut[3]  (.D(\shftOut_14[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft28_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_14[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft28_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_14[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft28_w[1]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_14_0_a2[7]  (.A(shft27_w[7]), 
        .B(fb_w_3), .C(N_566), .D(N_565), .Y(\shftOut_14[7] ));
    SLE \shftOut[0]  (.D(\shftOut_14[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft28_w[0]));
    CFG3 #( .INIT(8'h96) )  \shftOut_14_0_a2[5]  (.A(shft27_w[5]), .B(
        fb_w_7), .C(fb_w_1), .Y(\shftOut_14[5] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_171s_8s_0(
       Bit_Count_16dec_i_1,
       shft18_w,
       shft17_w,
       fb_w_1,
       fb_w_7,
       fb_w_3,
       fb_w_5,
       fb_w_0,
       fb_w_6,
       RSControl_0_NGRST,
       N_583,
       N_566,
       N_569,
       N_568,
       N_572,
       N_565,
       N_567,
       N_574
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft18_w;
input  [7:0] shft17_w;
input  fb_w_1;
input  fb_w_7;
input  fb_w_3;
input  fb_w_5;
input  fb_w_0;
input  fb_w_6;
input  RSControl_0_NGRST;
input  N_583;
input  N_566;
input  N_569;
input  N_568;
input  N_572;
input  N_565;
input  N_567;
input  N_574;

    wire VCC_net_1, \shftOut_41[3] , GND_net_1, \shftOut_41[4] , 
        \shftOut_41[5] , \shftOut_41[6] , \shftOut_41[7] , 
        \shftOut_41[0] , \shftOut_41[1] , \shftOut_41[2] ;
    
    CFG3 #( .INIT(8'h96) )  \shftOut_41_0_a2[2]  (.A(shft17_w[2]), .B(
        N_572), .C(N_565), .Y(\shftOut_41[2] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_41_0_a2[3]  (.A(shft17_w[3]), .B(
        N_583), .C(N_568), .Y(\shftOut_41[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_41_0_a2[0]  (.A(shft17_w[0]), .B(
        N_574), .C(N_569), .Y(\shftOut_41[0] ));
    SLE \shftOut[5]  (.D(\shftOut_41[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft18_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_41[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft18_w[6]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_41_0_a2[7]  (.A(shft17_w[7]), 
        .B(fb_w_1), .C(N_583), .D(N_566), .Y(\shftOut_41[7] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_41_0_a2[4]  (.A(shft17_w[4]), 
        .B(fb_w_7), .C(fb_w_1), .D(N_566), .Y(\shftOut_41[4] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_41[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft18_w[4]));
    CFG2 #( .INIT(4'h6) )  \shftOut_41_0_a2[5]  (.A(N_569), .B(
        shft17_w[5]), .Y(\shftOut_41[5] ));
    SLE \shftOut[7]  (.D(\shftOut_41[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft18_w[7]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_41_0_a2[1]  (.A(fb_w_3), .B(
        fb_w_5), .C(shft17_w[1]), .D(fb_w_0), .Y(\shftOut_41[1] ));
    SLE \shftOut[3]  (.D(\shftOut_41[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft18_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_41[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft18_w[2]));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h96) )  \shftOut_41_0_a2[6]  (.A(shft17_w[6]), .B(
        fb_w_6), .C(N_567), .Y(\shftOut_41[6] ));
    SLE \shftOut[1]  (.D(\shftOut_41[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft18_w[1]));
    SLE \shftOut[0]  (.D(\shftOut_41[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft18_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_97s_8s(
       Bit_Count_16dec_i_1,
       shft8_w,
       shft7_w,
       fb_w,
       RSControl_0_NGRST,
       N_564,
       N_567
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft8_w;
input  [7:0] shft7_w;
input  [7:0] fb_w;
input  RSControl_0_NGRST;
input  N_564;
input  N_567;

    wire VCC_net_1, \shftOut_26[3] , GND_net_1, \shftOut_26[4] , 
        \shftOut_26[5] , \shftOut_26[6] , \shftOut_26[7] , 
        \shftOut_26[0] , \shftOut_26[1] , \shftOut_26[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_26[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft8_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_26[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft8_w[6]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_26_0_a2[5]  (.A(fb_w[7]), .B(
        fb_w[6]), .C(shft7_w[5]), .D(fb_w[0]), .Y(\shftOut_26[5] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_26[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft8_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_26_0_a2[3]  (.A(fb_w[5]), .B(
        shft7_w[3]), .C(fb_w[4]), .Y(\shftOut_26[3] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_26_0_a2[0]  (.A(N_564), .B(
        shft7_w[0]), .Y(\shftOut_26[0] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_26_0_a2[1]  (.A(shft7_w[1]), .B(
        fb_w[2]), .C(N_567), .Y(\shftOut_26[1] ));
    SLE \shftOut[7]  (.D(\shftOut_26[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft8_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_26[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft8_w[3]));
    CFG3 #( .INIT(8'h96) )  \shftOut_26_0_a2[4]  (.A(shft7_w[4]), .B(
        fb_w[6]), .C(fb_w[5]), .Y(\shftOut_26[4] ));
    SLE \shftOut[2]  (.D(\shftOut_26[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft8_w[2]));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h6996) )  \shftOut_26_0_a2[6]  (.A(fb_w[7]), .B(
        fb_w[1]), .C(shft7_w[6]), .D(fb_w[0]), .Y(\shftOut_26[6] ));
    SLE \shftOut[1]  (.D(\shftOut_26[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft8_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_26_0_a2[2]  (.A(shft7_w[2]), .B(
        fb_w[4]), .C(fb_w[3]), .Y(\shftOut_26[2] ));
    SLE \shftOut[0]  (.D(\shftOut_26[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft8_w[0]));
    CFG2 #( .INIT(4'h6) )  \shftOut_26_0_a2[7]  (.A(fb_w[1]), .B(
        shft7_w[7]), .Y(\shftOut_26[7] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_235s_8s_0(
       Bit_Count_16dec_i_1,
       shft25_w,
       shft24_w,
       fb_w_1,
       fb_w_6,
       fb_w_7,
       fb_w_0,
       fb_w_3,
       fb_w_5,
       fb_w_4,
       RSControl_0_NGRST,
       N_564,
       N_567
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft25_w;
input  [7:0] shft24_w;
input  fb_w_1;
input  fb_w_6;
input  fb_w_7;
input  fb_w_0;
input  fb_w_3;
input  fb_w_5;
input  fb_w_4;
input  RSControl_0_NGRST;
input  N_564;
input  N_567;

    wire VCC_net_1, \shftOut_23[3] , GND_net_1, \shftOut_23[4] , 
        \shftOut_23[5] , \shftOut_23[6] , \shftOut_23[7] , 
        \shftOut_23[0] , \shftOut_23[1] , \shftOut_23[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_23[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft25_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_23[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft25_w[6]));
    CFG2 #( .INIT(4'h6) )  \shftOut_23_0_a2[5]  (.A(N_564), .B(
        shft24_w[5]), .Y(\shftOut_23[5] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_23[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft25_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_23_0_a2[3]  (.A(fb_w_7), .B(
        shft24_w[3]), .C(fb_w_0), .Y(\shftOut_23[3] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_23_0_a2[0]  (.A(shft24_w[0]), 
        .B(fb_w_4), .C(fb_w_0), .D(N_567), .Y(\shftOut_23[0] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_23_0_a2[1]  (.A(shft24_w[1]), 
        .B(fb_w_3), .C(fb_w_5), .D(N_564), .Y(\shftOut_23[1] ));
    SLE \shftOut[7]  (.D(\shftOut_23[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft25_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_23[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft25_w[3]));
    CFG2 #( .INIT(4'h6) )  \shftOut_23_0_a2[4]  (.A(fb_w_1), .B(
        shft24_w[4]), .Y(\shftOut_23[4] ));
    SLE \shftOut[2]  (.D(\shftOut_23[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft25_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_23[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft25_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_23_0_a2[6]  (.A(shft24_w[6]), .B(
        fb_w_0), .C(N_567), .Y(\shftOut_23[6] ));
    SLE \shftOut[0]  (.D(\shftOut_23[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft25_w[0]));
    CFG2 #( .INIT(4'h6) )  \shftOut_23_0_a2[2]  (.A(fb_w_6), .B(
        shft24_w[2]), .Y(\shftOut_23[2] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_23_0_a2[7]  (.A(shft24_w[7]), .B(
        fb_w_3), .C(N_564), .Y(\shftOut_23[7] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_32s_8s(
       Bit_Count_16dec_i_1,
       shft15_w,
       shft14_w,
       fb_w_3,
       fb_w_6,
       fb_w_0,
       fb_w_7,
       fb_w_1,
       fb_w_2,
       RSControl_0_NGRST,
       N_566,
       N_565,
       N_568,
       N_573
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft15_w;
input  [7:0] shft14_w;
input  fb_w_3;
input  fb_w_6;
input  fb_w_0;
input  fb_w_7;
input  fb_w_1;
input  fb_w_2;
input  RSControl_0_NGRST;
input  N_566;
input  N_565;
input  N_568;
input  N_573;

    wire VCC_net_1, \shftOut_44[3] , GND_net_1, \shftOut_44[4] , 
        \shftOut_44[5] , \shftOut_44[6] , \shftOut_44[7] , 
        \shftOut_44[0] , \shftOut_44[1] , \shftOut_44[2] ;
    
    CFG2 #( .INIT(4'h6) )  \shftOut_44_0_a2[1]  (.A(fb_w_3), .B(
        shft14_w[1]), .Y(\shftOut_44[1] ));
    SLE \shftOut[5]  (.D(\shftOut_44[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft15_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_44[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft15_w[6]));
    CFG3 #( .INIT(8'h96) )  \shftOut_44_0_a2[6]  (.A(shft14_w[6]), .B(
        fb_w_7), .C(fb_w_1), .Y(\shftOut_44[6] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_44[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft15_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_44_0_a2[2]  (.A(shft14_w[2]), .B(
        N_568), .C(N_565), .Y(\shftOut_44[2] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_44_0_a2[3]  (.A(shft14_w[3]), .B(
        fb_w_7), .C(N_566), .Y(\shftOut_44[3] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_44_0_a2[0]  (.A(shft14_w[0]), 
        .B(fb_w_3), .C(N_566), .D(N_565), .Y(\shftOut_44[0] ));
    SLE \shftOut[7]  (.D(\shftOut_44[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft15_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_44[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft15_w[3]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_44_0_a2[7]  (.A(shft14_w[7]), 
        .B(fb_w_2), .C(fb_w_3), .D(N_573), .Y(\shftOut_44[7] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_44_0_a2[4]  (.A(N_565), .B(
        shft14_w[4]), .Y(\shftOut_44[4] ));
    SLE \shftOut[2]  (.D(\shftOut_44[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft15_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_44[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft15_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_44_0_a2[5]  (.A(fb_w_6), .B(
        shft14_w[5]), .C(fb_w_0), .Y(\shftOut_44[5] ));
    SLE \shftOut[0]  (.D(\shftOut_44[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft15_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_165s_8s_0(
       Bit_Count_16dec_i_1,
       shft23_w,
       shft22_w,
       fb_w,
       RSControl_0_NGRST,
       N_574,
       N_566,
       N_568,
       N_564,
       N_570,
       N_567,
       N_565,
       N_588
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft23_w;
input  [7:0] shft22_w;
input  [7:0] fb_w;
input  RSControl_0_NGRST;
output N_574;
input  N_566;
input  N_568;
input  N_564;
input  N_570;
input  N_567;
input  N_565;
input  N_588;

    wire VCC_net_1, \shftOut_29[3] , GND_net_1, \shftOut_29[4] , 
        \shftOut_29[5] , \shftOut_29[6] , \shftOut_29[7] , 
        \shftOut_29[0] , \shftOut_29[1] , \shftOut_29[2] ;
    
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[5]  (.A(shft22_w[5]), 
        .B(fb_w[4]), .C(N_588), .D(N_565), .Y(\shftOut_29[5] ));
    SLE \shftOut[5]  (.D(\shftOut_29[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft23_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_29[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft23_w[6]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[3]  (.A(fb_w[2]), .B(
        shft22_w[3]), .C(N_567), .D(N_565), .Y(\shftOut_29[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_29_0_a2[0]  (.A(shft22_w[0]), .B(
        N_574), .C(N_564), .Y(\shftOut_29[0] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_29[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft23_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_29_0_a2[1]  (.A(shft22_w[1]), .B(
        fb_w[7]), .C(N_568), .Y(\shftOut_29[1] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_29_0_a2_0[0]  (.A(fb_w[6]), .B(
        fb_w[1]), .Y(N_574));
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[4]  (.A(shft22_w[4]), 
        .B(fb_w[2]), .C(fb_w[3]), .D(N_566), .Y(\shftOut_29[4] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[6]  (.A(shft22_w[6]), 
        .B(fb_w[1]), .C(fb_w[5]), .D(N_566), .Y(\shftOut_29[6] ));
    SLE \shftOut[7]  (.D(\shftOut_29[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft23_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_29[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft23_w[3]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[2]  (.A(shft22_w[2]), 
        .B(fb_w[7]), .C(fb_w[1]), .D(N_570), .Y(\shftOut_29[2] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_29_0_a2[7]  (.A(shft22_w[7]), 
        .B(fb_w[0]), .C(fb_w[1]), .D(N_565), .Y(\shftOut_29[7] ));
    SLE \shftOut[2]  (.D(\shftOut_29[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft23_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_29[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft23_w[1]));
    SLE \shftOut[0]  (.D(\shftOut_29[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft23_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_13s_8s_0(
       Bit_Count_16dec_i_1,
       shft26_w,
       fb_w,
       shft25_w,
       RSControl_0_NGRST,
       N_576,
       N_583,
       N_574,
       N_572,
       N_566,
       N_575,
       N_569
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft26_w;
input  [7:0] fb_w;
input  [7:0] shft25_w;
input  RSControl_0_NGRST;
output N_576;
output N_583;
input  N_574;
input  N_572;
input  N_566;
input  N_575;
input  N_569;

    wire VCC_net_1, \shftOut_20[3] , GND_net_1, \shftOut_20[4] , 
        \shftOut_20[5] , \shftOut_20[6] , \shftOut_20[7] , 
        \shftOut_20[0] , \shftOut_20[1] , \shftOut_20[2] ;
    
    CFG2 #( .INIT(4'h6) )  \shftOut_20_0_a2[0]  (.A(N_583), .B(
        shft25_w[0]), .Y(\shftOut_20[0] ));
    SLE \shftOut[5]  (.D(\shftOut_20[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft26_w[5]));
    CFG3 #( .INIT(8'h96) )  \shftOut_20_0_a2[1]  (.A(shft25_w[1]), .B(
        fb_w[5]), .C(N_574), .Y(\shftOut_20[1] ));
    SLE \shftOut[6]  (.D(\shftOut_20[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft26_w[6]));
    CFG2 #( .INIT(4'h6) )  \shftOut_20_0_a2_0[0]  (.A(fb_w[5]), .B(
        fb_w[0]), .Y(N_583));
    CFG4 #( .INIT(16'h6996) )  \shftOut_20_0_a2[4]  (.A(shft25_w[4]), 
        .B(fb_w[7]), .C(fb_w[1]), .D(N_572), .Y(\shftOut_20[4] ));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h6) )  \shftOut_20_0_a2_0[7]  (.A(fb_w[7]), .B(
        fb_w[4]), .Y(N_576));
    SLE \shftOut[4]  (.D(\shftOut_20[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft26_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_20_0_a2[6]  (.A(shft25_w[6]), .B(
        fb_w[3]), .C(N_566), .Y(\shftOut_20[6] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_20_0_a2[2]  (.A(shft25_w[2]), .B(
        fb_w[6]), .C(N_569), .Y(\shftOut_20[2] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_20_0_a2[7]  (.A(N_576), .B(
        shft25_w[7]), .Y(\shftOut_20[7] ));
    SLE \shftOut[7]  (.D(\shftOut_20[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft26_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_20[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft26_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_20[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft26_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_20[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft26_w[1]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_20_0_a2[5]  (.A(fb_w[3]), .B(
        fb_w[5]), .C(shft25_w[5]), .D(fb_w[2]), .Y(\shftOut_20[5] ));
    SLE \shftOut[0]  (.D(\shftOut_20[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft26_w[0]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_20_0_a2[3]  (.A(shft25_w[3]), 
        .B(fb_w[0]), .C(fb_w[6]), .D(N_575), .Y(\shftOut_20[3] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_86s_8s_0(
       Bit_Count_16dec_i_1,
       shft13_w,
       shft12_w,
       fb_w,
       RSControl_0_NGRST,
       N_568,
       N_567,
       N_574,
       N_569,
       N_576,
       N_564,
       N_565,
       N_570,
       N_575
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft13_w;
input  [7:0] shft12_w;
input  [7:1] fb_w;
input  RSControl_0_NGRST;
input  N_568;
input  N_567;
input  N_574;
input  N_569;
input  N_576;
input  N_564;
input  N_565;
input  N_570;
input  N_575;

    wire VCC_net_1, \shftOut_11[3] , GND_net_1, \shftOut_11[4] , 
        \shftOut_11[5] , \shftOut_11[6] , \shftOut_11[7] , 
        \shftOut_11[0] , \shftOut_11[1] , \shftOut_11[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_11[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft13_w[5]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[3]  (.A(shft12_w[3]), 
        .B(fb_w[2]), .C(fb_w[6]), .D(N_575), .Y(\shftOut_11[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[2]  (.A(shft12_w[2]), .B(
        N_574), .C(N_569), .Y(\shftOut_11[2] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[6]  (.A(shft12_w[6]), .B(
        fb_w[5]), .C(N_570), .Y(\shftOut_11[6] ));
    SLE \shftOut[6]  (.D(\shftOut_11[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft13_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_11[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft13_w[4]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[7]  (.A(shft12_w[7]), 
        .B(fb_w[2]), .C(fb_w[1]), .D(N_565), .Y(\shftOut_11[7] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[5]  (.A(shft12_w[5]), 
        .B(fb_w[4]), .C(fb_w[5]), .D(N_567), .Y(\shftOut_11[5] ));
    SLE \shftOut[7]  (.D(\shftOut_11[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft13_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_11[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft13_w[3]));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[1]  (.A(shft12_w[1]), .B(
        fb_w[7]), .C(N_570), .Y(\shftOut_11[1] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_11_0_a2[0]  (.A(shft12_w[0]), .B(
        fb_w[2]), .C(N_568), .Y(\shftOut_11[0] ));
    SLE \shftOut[2]  (.D(\shftOut_11[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft13_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_11[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft13_w[1]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_11_0_a2[4]  (.A(shft12_w[4]), 
        .B(fb_w[3]), .C(N_576), .D(N_564), .Y(\shftOut_11[4] ));
    SLE \shftOut[0]  (.D(\shftOut_11[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft13_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_113s_8s(
       Bit_Count_16dec_i_1,
       shft16_w,
       shft15_w,
       fb_w_0,
       fb_w_7,
       fb_w_1,
       RSControl_0_NGRST,
       N_566,
       N_567,
       N_565,
       N_574,
       N_576,
       N_583,
       N_569,
       N_564,
       N_572,
       N_568
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft16_w;
input  [7:0] shft15_w;
input  fb_w_0;
input  fb_w_7;
input  fb_w_1;
input  RSControl_0_NGRST;
input  N_566;
input  N_567;
input  N_565;
input  N_574;
input  N_576;
input  N_583;
input  N_569;
input  N_564;
input  N_572;
input  N_568;

    wire VCC_net_1, \shftOut_47[3] , GND_net_1, \shftOut_47[4] , 
        \shftOut_47[5] , \shftOut_47[6] , \shftOut_47[7] , 
        \shftOut_47[0] , \shftOut_47[1] , \shftOut_47[2] ;
    
    CFG4 #( .INIT(16'h6996) )  \shftOut_47_0_a2[7]  (.A(N_566), .B(
        shft15_w[7]), .C(N_567), .D(N_565), .Y(\shftOut_47[7] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_47_0_a2[4]  (.A(N_583), .B(
        shft15_w[4]), .Y(\shftOut_47[4] ));
    SLE \shftOut[5]  (.D(\shftOut_47[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft16_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_47[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft16_w[6]));
    CFG3 #( .INIT(8'h96) )  \shftOut_47_0_a2[5]  (.A(shft15_w[5]), .B(
        fb_w_0), .C(N_574), .Y(\shftOut_47[5] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_47[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft16_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_47_0_a2[1]  (.A(shft15_w[1]), .B(
        N_572), .C(N_567), .Y(\shftOut_47[1] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_47_0_a2[6]  (.A(shft15_w[6]), 
        .B(fb_w_7), .C(fb_w_1), .D(N_564), .Y(\shftOut_47[6] ));
    SLE \shftOut[7]  (.D(\shftOut_47[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft16_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_47[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft16_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_47[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft16_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_47[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft16_w[1]));
    SLE \shftOut[0]  (.D(\shftOut_47[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft16_w[0]));
    CFG3 #( .INIT(8'h96) )  \shftOut_47_0_a2[2]  (.A(shft15_w[2]), .B(
        fb_w_7), .C(N_568), .Y(\shftOut_47[2] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_47_0_a2[3]  (.A(N_576), .B(
        shft15_w[3]), .Y(\shftOut_47[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_47_0_a2[0]  (.A(N_569), .B(
        shft15_w[0]), .C(N_566), .Y(\shftOut_47[0] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_42s_8s_0(
       Bit_Count_16dec_i_1,
       shft21_w,
       shft20_w,
       fb_w_1,
       fb_w_3,
       fb_w_5,
       fb_w_0,
       fb_w_4,
       RSControl_0_NGRST,
       N_576,
       N_564,
       N_567,
       N_565,
       N_588,
       N_570,
       N_568,
       N_575
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft21_w;
input  [7:0] shft20_w;
input  fb_w_1;
input  fb_w_3;
input  fb_w_5;
input  fb_w_0;
input  fb_w_4;
input  RSControl_0_NGRST;
input  N_576;
input  N_564;
input  N_567;
input  N_565;
input  N_588;
input  N_570;
input  N_568;
input  N_575;

    wire VCC_net_1, \shftOut_35[3] , GND_net_1, \shftOut_35[4] , 
        \shftOut_35[5] , \shftOut_35[6] , \shftOut_35[7] , 
        \shftOut_35[0] , \shftOut_35[1] , \shftOut_35[2] ;
    
    CFG4 #( .INIT(16'h6996) )  \shftOut_35_0_a2[7]  (.A(shft20_w[7]), 
        .B(fb_w_5), .C(fb_w_0), .D(N_568), .Y(\shftOut_35[7] ));
    SLE \shftOut[5]  (.D(\shftOut_35[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft21_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_35[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft21_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_35[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft21_w[4]));
    CFG2 #( .INIT(4'h6) )  \shftOut_35_0_a2[5]  (.A(N_570), .B(
        shft20_w[5]), .Y(\shftOut_35[5] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[4]  (.A(shft20_w[4]), .B(
        fb_w_3), .C(N_567), .Y(\shftOut_35[4] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[3]  (.A(shft20_w[3]), .B(
        N_576), .C(N_564), .Y(\shftOut_35[3] ));
    SLE \shftOut[7]  (.D(\shftOut_35[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft21_w[7]));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[6]  (.A(N_567), .B(
        shft20_w[6]), .C(N_565), .Y(\shftOut_35[6] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[2]  (.A(shft20_w[2]), .B(
        fb_w_4), .C(N_575), .Y(\shftOut_35[2] ));
    SLE \shftOut[3]  (.D(\shftOut_35[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft21_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_35[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft21_w[2]));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[0]  (.A(shft20_w[0]), .B(
        fb_w_1), .C(N_576), .Y(\shftOut_35[0] ));
    SLE \shftOut[1]  (.D(\shftOut_35[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft21_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[1]  (.A(shft20_w[1]), .B(
        N_588), .C(N_565), .Y(\shftOut_35[1] ));
    SLE \shftOut[0]  (.D(\shftOut_35[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft21_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_42s_8s(
       Bit_Count_16dec_i_1,
       shft11_w,
       shft10_w,
       fb_w_1,
       fb_w_3,
       fb_w_5,
       fb_w_0,
       fb_w_4,
       RSControl_0_NGRST,
       N_576,
       N_564,
       N_567,
       N_565,
       N_588,
       N_570,
       N_568,
       N_575
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft11_w;
input  [7:0] shft10_w;
input  fb_w_1;
input  fb_w_3;
input  fb_w_5;
input  fb_w_0;
input  fb_w_4;
input  RSControl_0_NGRST;
input  N_576;
input  N_564;
input  N_567;
input  N_565;
input  N_588;
input  N_570;
input  N_568;
input  N_575;

    wire VCC_net_1, \shftOut_35[3] , GND_net_1, \shftOut_35[4] , 
        \shftOut_35[5] , \shftOut_35[6] , \shftOut_35[7] , 
        \shftOut_35[0] , \shftOut_35[1] , \shftOut_35[2] ;
    
    CFG4 #( .INIT(16'h6996) )  \shftOut_35_0_a2[7]  (.A(shft10_w[7]), 
        .B(fb_w_5), .C(fb_w_0), .D(N_568), .Y(\shftOut_35[7] ));
    SLE \shftOut[5]  (.D(\shftOut_35[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft11_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_35[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft11_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_35[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft11_w[4]));
    CFG2 #( .INIT(4'h6) )  \shftOut_35_0_a2[5]  (.A(N_570), .B(
        shft10_w[5]), .Y(\shftOut_35[5] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[4]  (.A(shft10_w[4]), .B(
        fb_w_3), .C(N_567), .Y(\shftOut_35[4] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[3]  (.A(shft10_w[3]), .B(
        N_576), .C(N_564), .Y(\shftOut_35[3] ));
    SLE \shftOut[7]  (.D(\shftOut_35[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft11_w[7]));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[6]  (.A(N_567), .B(
        shft10_w[6]), .C(N_565), .Y(\shftOut_35[6] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[2]  (.A(shft10_w[2]), .B(
        fb_w_4), .C(N_575), .Y(\shftOut_35[2] ));
    SLE \shftOut[3]  (.D(\shftOut_35[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft11_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_35[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft11_w[2]));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[0]  (.A(shft10_w[0]), .B(
        fb_w_1), .C(N_576), .Y(\shftOut_35[0] ));
    SLE \shftOut[1]  (.D(\shftOut_35[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft11_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_35_0_a2[1]  (.A(shft10_w[1]), .B(
        N_588), .C(N_565), .Y(\shftOut_35[1] ));
    SLE \shftOut[0]  (.D(\shftOut_35[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft11_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_127s_8s_0(
       Bit_Count_16dec_i_1,
       shft30_w,
       shft29_w,
       dInp_reg_w_3,
       dInp_reg_w_2,
       dInp_reg_w_0,
       pre_fb_w_3,
       pre_fb_w_2,
       pre_fb_w_0,
       fb_w_4,
       fb_w_7,
       fb_w_1,
       fb_w_5,
       fb_w_0,
       RSControl_0_NGRST,
       N_564,
       N_570,
       N_565,
       N_567,
       N_566,
       N_569
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft30_w;
input  [7:0] shft29_w;
input  dInp_reg_w_3;
input  dInp_reg_w_2;
input  dInp_reg_w_0;
input  pre_fb_w_3;
input  pre_fb_w_2;
input  pre_fb_w_0;
input  fb_w_4;
input  fb_w_7;
input  fb_w_1;
input  fb_w_5;
input  fb_w_0;
input  RSControl_0_NGRST;
input  N_564;
output N_570;
output N_565;
output N_567;
output N_566;
input  N_569;

    wire VCC_net_1, \shftOut_8[3] , GND_net_1, \shftOut_8[4] , 
        \shftOut_8[5] , \shftOut_8[6] , \shftOut_8[7] , \shftOut_8[0] , 
        \shftOut_8[1] , \shftOut_8[2] ;
    
    CFG4 #( .INIT(16'h6996) )  \shftOut_8_0_a2_1[5]  (.A(fb_w_4), .B(
        N_564), .C(pre_fb_w_3), .D(dInp_reg_w_3), .Y(N_570));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2_0[5]  (.A(dInp_reg_w_0), 
        .B(fb_w_1), .C(pre_fb_w_0), .Y(N_567));
    SLE \shftOut[5]  (.D(\shftOut_8[5] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft30_w[5]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_8_0_a2[1]  (.A(N_567), .B(
        N_569), .C(shft29_w[1]), .D(N_566), .Y(\shftOut_8[1] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2[5]  (.A(N_570), .B(
        shft29_w[5]), .C(N_567), .Y(\shftOut_8[5] ));
    SLE \shftOut[6]  (.D(\shftOut_8[6] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft30_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_8[4] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft30_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2_0[1]  (.A(dInp_reg_w_3), 
        .B(fb_w_4), .C(pre_fb_w_3), .Y(N_566));
    SLE \shftOut[7]  (.D(\shftOut_8[7] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft30_w[7]));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2[7]  (.A(shft29_w[7]), .B(
        fb_w_5), .C(N_567), .Y(\shftOut_8[7] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_8_0_a2[0]  (.A(N_570), .B(
        shft29_w[0]), .Y(\shftOut_8[0] ));
    SLE \shftOut[3]  (.D(\shftOut_8[3] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft30_w[3]));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2_0[2]  (.A(dInp_reg_w_2), 
        .B(fb_w_7), .C(pre_fb_w_2), .Y(N_565));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2[4]  (.A(N_569), .B(
        shft29_w[4]), .C(N_567), .Y(\shftOut_8[4] ));
    SLE \shftOut[2]  (.D(\shftOut_8[2] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft30_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_8[1] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft30_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2[3]  (.A(shft29_w[3]), .B(
        fb_w_1), .C(N_570), .Y(\shftOut_8[3] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_8_0_a2[2]  (.A(fb_w_0), .B(
        shft29_w[2]), .C(N_567), .D(N_565), .Y(\shftOut_8[2] ));
    SLE \shftOut[0]  (.D(\shftOut_8[0] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft30_w[0]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_8_0_a2[6]  (.A(fb_w_4), .B(
        shft29_w[6]), .C(N_569), .D(N_567), .Y(\shftOut_8[6] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_97s_8s_0(
       Bit_Count_16dec_i_1,
       shft24_w,
       shft23_w,
       fb_w,
       RSControl_0_NGRST,
       N_564,
       N_567
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft24_w;
input  [7:0] shft23_w;
input  [7:0] fb_w;
input  RSControl_0_NGRST;
input  N_564;
input  N_567;

    wire VCC_net_1, \shftOut_26[3] , GND_net_1, \shftOut_26[4] , 
        \shftOut_26[5] , \shftOut_26[6] , \shftOut_26[7] , 
        \shftOut_26[0] , \shftOut_26[1] , \shftOut_26[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_26[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft24_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_26[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft24_w[6]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_26_0_a2[5]  (.A(fb_w[7]), .B(
        fb_w[6]), .C(shft23_w[5]), .D(fb_w[0]), .Y(\shftOut_26[5] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_26[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft24_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_26_0_a2[3]  (.A(fb_w[5]), .B(
        shft23_w[3]), .C(fb_w[4]), .Y(\shftOut_26[3] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_26_0_a2[0]  (.A(N_564), .B(
        shft23_w[0]), .Y(\shftOut_26[0] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_26_0_a2[1]  (.A(shft23_w[1]), .B(
        fb_w[2]), .C(N_567), .Y(\shftOut_26[1] ));
    SLE \shftOut[7]  (.D(\shftOut_26[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft24_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_26[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft24_w[3]));
    CFG3 #( .INIT(8'h96) )  \shftOut_26_0_a2[4]  (.A(shft23_w[4]), .B(
        fb_w[6]), .C(fb_w[5]), .Y(\shftOut_26[4] ));
    SLE \shftOut[2]  (.D(\shftOut_26[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft24_w[2]));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h6996) )  \shftOut_26_0_a2[6]  (.A(fb_w[7]), .B(
        fb_w[1]), .C(shft23_w[6]), .D(fb_w[0]), .Y(\shftOut_26[6] ));
    SLE \shftOut[1]  (.D(\shftOut_26[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft24_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_26_0_a2[2]  (.A(shft23_w[2]), .B(
        fb_w[4]), .C(fb_w[3]), .Y(\shftOut_26[2] ));
    SLE \shftOut[0]  (.D(\shftOut_26[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft24_w[0]));
    CFG2 #( .INIT(4'h6) )  \shftOut_26_0_a2[7]  (.A(fb_w[1]), .B(
        shft23_w[7]), .Y(\shftOut_26[7] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_171s_8s(
       Bit_Count_16dec_i_1,
       shft14_w,
       shft13_w,
       fb_w_1,
       fb_w_7,
       fb_w_3,
       fb_w_5,
       fb_w_0,
       fb_w_6,
       RSControl_0_NGRST,
       N_583,
       N_566,
       N_569,
       N_568,
       N_572,
       N_565,
       N_567,
       N_574
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft14_w;
input  [7:0] shft13_w;
input  fb_w_1;
input  fb_w_7;
input  fb_w_3;
input  fb_w_5;
input  fb_w_0;
input  fb_w_6;
input  RSControl_0_NGRST;
input  N_583;
input  N_566;
input  N_569;
input  N_568;
input  N_572;
input  N_565;
input  N_567;
input  N_574;

    wire VCC_net_1, \shftOut_41[3] , GND_net_1, \shftOut_41[4] , 
        \shftOut_41[5] , \shftOut_41[6] , \shftOut_41[7] , 
        \shftOut_41[0] , \shftOut_41[1] , \shftOut_41[2] ;
    
    CFG3 #( .INIT(8'h96) )  \shftOut_41_0_a2[2]  (.A(shft13_w[2]), .B(
        N_572), .C(N_565), .Y(\shftOut_41[2] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_41_0_a2[3]  (.A(shft13_w[3]), .B(
        N_583), .C(N_568), .Y(\shftOut_41[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_41_0_a2[0]  (.A(shft13_w[0]), .B(
        N_574), .C(N_569), .Y(\shftOut_41[0] ));
    SLE \shftOut[5]  (.D(\shftOut_41[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft14_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_41[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft14_w[6]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_41_0_a2[7]  (.A(shft13_w[7]), 
        .B(fb_w_1), .C(N_583), .D(N_566), .Y(\shftOut_41[7] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_41_0_a2[4]  (.A(shft13_w[4]), 
        .B(fb_w_7), .C(fb_w_1), .D(N_566), .Y(\shftOut_41[4] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_41[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft14_w[4]));
    CFG2 #( .INIT(4'h6) )  \shftOut_41_0_a2[5]  (.A(N_569), .B(
        shft13_w[5]), .Y(\shftOut_41[5] ));
    SLE \shftOut[7]  (.D(\shftOut_41[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft14_w[7]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_41_0_a2[1]  (.A(fb_w_3), .B(
        fb_w_5), .C(shft13_w[1]), .D(fb_w_0), .Y(\shftOut_41[1] ));
    SLE \shftOut[3]  (.D(\shftOut_41[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft14_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_41[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft14_w[2]));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h96) )  \shftOut_41_0_a2[6]  (.A(shft13_w[6]), .B(
        fb_w_6), .C(N_567), .Y(\shftOut_41[6] ));
    SLE \shftOut[1]  (.D(\shftOut_41[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft14_w[1]));
    SLE \shftOut[0]  (.D(\shftOut_41[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft14_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_8s_8s_0(
       Bit_Count_16dec_i_1,
       shft22_w,
       shft21_w,
       fb_w_2,
       fb_w_5,
       fb_w_3,
       fb_w_6,
       fb_w_0,
       fb_w_7,
       fb_w_1,
       RSControl_0_NGRST,
       N_566,
       N_565
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft22_w;
input  [7:0] shft21_w;
input  fb_w_2;
input  fb_w_5;
input  fb_w_3;
input  fb_w_6;
input  fb_w_0;
input  fb_w_7;
input  fb_w_1;
input  RSControl_0_NGRST;
input  N_566;
input  N_565;

    wire VCC_net_1, \shftOut_32[3] , GND_net_1, \shftOut_32[4] , 
        \shftOut_32[5] , \shftOut_32[6] , \shftOut_32[7] , 
        \shftOut_32[0] , \shftOut_32[1] , \shftOut_32[2] ;
    
    CFG3 #( .INIT(8'h96) )  \shftOut_32_0_a2[0]  (.A(shft21_w[0]), .B(
        fb_w_6), .C(N_565), .Y(\shftOut_32[0] ));
    SLE \shftOut[5]  (.D(\shftOut_32[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft22_w[5]));
    CFG2 #( .INIT(4'h6) )  \shftOut_32_0_a2[1]  (.A(fb_w_5), .B(
        shft21_w[1]), .Y(\shftOut_32[1] ));
    SLE \shftOut[6]  (.D(\shftOut_32[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft22_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_32[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft22_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_32_0_a2[7]  (.A(shft21_w[7]), .B(
        N_566), .C(N_565), .Y(\shftOut_32[7] ));
    SLE \shftOut[7]  (.D(\shftOut_32[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft22_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_32[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft22_w[3]));
    CFG2 #( .INIT(4'h6) )  \shftOut_32_0_a2[5]  (.A(fb_w_2), .B(
        shft21_w[5]), .Y(\shftOut_32[5] ));
    SLE \shftOut[2]  (.D(\shftOut_32[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft22_w[2]));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h96) )  \shftOut_32_0_a2[4]  (.A(shft21_w[4]), .B(
        fb_w_7), .C(fb_w_1), .Y(\shftOut_32[4] ));
    SLE \shftOut[1]  (.D(\shftOut_32[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft22_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_32_0_a2[3]  (.A(fb_w_6), .B(
        shft21_w[3]), .C(fb_w_0), .Y(\shftOut_32[3] ));
    SLE \shftOut[0]  (.D(\shftOut_32[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft22_w[0]));
    CFG2 #( .INIT(4'h6) )  \shftOut_32_0_a2[6]  (.A(fb_w_3), .B(
        shft21_w[6]), .Y(\shftOut_32[6] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_32_0_a2[2]  (.A(N_565), .B(
        shft21_w[2]), .Y(\shftOut_32[2] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_54s_8s(
       Bit_Count_16dec_i_1,
       shft12_w,
       shft11_w,
       fb_w_5,
       fb_w_2,
       fb_w_0,
       fb_w_1,
       fb_w_7,
       RSControl_0_NGRST,
       N_568,
       N_575,
       N_566,
       N_573,
       N_567,
       N_569,
       N_572,
       N_565,
       N_588
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft12_w;
input  [7:0] shft11_w;
input  fb_w_5;
input  fb_w_2;
input  fb_w_0;
input  fb_w_1;
input  fb_w_7;
input  RSControl_0_NGRST;
input  N_568;
input  N_575;
input  N_566;
input  N_573;
input  N_567;
input  N_569;
input  N_572;
input  N_565;
input  N_588;

    wire VCC_net_1, \shftOut_38[3] , GND_net_1, \shftOut_38[4] , 
        \shftOut_38[5] , \shftOut_38[6] , \shftOut_38[7] , 
        \shftOut_38[0] , \shftOut_38[1] , \shftOut_38[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_38[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft12_w[5]));
    CFG3 #( .INIT(8'h96) )  \shftOut_38_0_a2[7]  (.A(fb_w_5), .B(
        shft11_w[7]), .C(fb_w_2), .Y(\shftOut_38[7] ));
    SLE \shftOut[6]  (.D(\shftOut_38[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft12_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_38[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft12_w[4]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_38_0_a2[5]  (.A(shft11_w[5]), 
        .B(fb_w_0), .C(N_575), .D(N_566), .Y(\shftOut_38[5] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_38_0_a2[4]  (.A(N_569), .B(
        shft11_w[4]), .C(N_568), .Y(\shftOut_38[4] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_38_0_a2[3]  (.A(shft11_w[3]), 
        .B(fb_w_2), .C(fb_w_1), .D(N_573), .Y(\shftOut_38[3] ));
    SLE \shftOut[7]  (.D(\shftOut_38[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft12_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_38[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft12_w[3]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_38_0_a2[6]  (.A(shft11_w[6]), 
        .B(fb_w_1), .C(N_572), .D(N_565), .Y(\shftOut_38[6] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_38_0_a2[2]  (.A(fb_w_0), .B(
        shft11_w[2]), .C(N_573), .D(N_567), .Y(\shftOut_38[2] ));
    SLE \shftOut[2]  (.D(\shftOut_38[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft12_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_38[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft12_w[1]));
    CFG2 #( .INIT(4'h6) )  \shftOut_38_0_a2[0]  (.A(N_568), .B(
        shft11_w[0]), .Y(\shftOut_38[0] ));
    SLE \shftOut[0]  (.D(\shftOut_38[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft12_w[0]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_38_0_a2[1]  (.A(shft11_w[1]), 
        .B(fb_w_7), .C(N_588), .D(N_566), .Y(\shftOut_38[1] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_30s_8s(
       Bit_Count_16dec_i_1,
       shft5_w,
       shftOut_17_1,
       shft4_w,
       fb_w_0,
       fb_w_5,
       fb_w_3,
       fb_w_6,
       RSControl_0_NGRST,
       N_566,
       N_565,
       N_572,
       N_575,
       N_574,
       N_564
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft5_w;
input  [2:2] shftOut_17_1;
input  [7:0] shft4_w;
input  fb_w_0;
input  fb_w_5;
input  fb_w_3;
input  fb_w_6;
input  RSControl_0_NGRST;
input  N_566;
input  N_565;
input  N_572;
input  N_575;
input  N_574;
input  N_564;

    wire VCC_net_1, \shftOut_17[3] , GND_net_1, \shftOut_17[4] , 
        \shftOut_17[5] , \shftOut_17[6] , \shftOut_17[7] , 
        \shftOut_17[0] , \shftOut_17[1] , \shftOut_17[2] ;
    
    CFG4 #( .INIT(16'h6996) )  \shftOut_17_0_a2[6]  (.A(shft4_w[6]), 
        .B(fb_w_3), .C(fb_w_5), .D(N_572), .Y(\shftOut_17[6] ));
    SLE \shftOut[5]  (.D(\shftOut_17[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft5_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_17[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft5_w[6]));
    CFG3 #( .INIT(8'h96) )  \shftOut_17_0_a2[7]  (.A(fb_w_5), .B(
        shft4_w[7]), .C(fb_w_3), .Y(\shftOut_17[7] ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h96) )  \shftOut_17_0_a2[5]  (.A(N_575), .B(
        shft4_w[5]), .C(N_572), .Y(\shftOut_17[5] ));
    SLE \shftOut[4]  (.D(\shftOut_17[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft5_w[4]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_17_0_a2[1]  (.A(shft4_w[1]), 
        .B(fb_w_0), .C(N_566), .D(N_565), .Y(\shftOut_17[1] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_17_0_a2[0]  (.A(N_566), .B(
        shft4_w[0]), .Y(\shftOut_17[0] ));
    SLE \shftOut[7]  (.D(\shftOut_17[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft5_w[7]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_17_0_a2[4]  (.A(shft4_w[4]), 
        .B(fb_w_6), .C(N_575), .D(N_564), .Y(\shftOut_17[4] ));
    SLE \shftOut[3]  (.D(\shftOut_17[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft5_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_17[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft5_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_17[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft5_w[1]));
    SLE \shftOut[0]  (.D(\shftOut_17[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft5_w[0]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_17_0_a2[3]  (.A(shft4_w[3]), 
        .B(fb_w_5), .C(N_574), .D(N_564), .Y(\shftOut_17[3] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_17_0_a2[2]  (.A(shftOut_17_1[2]), 
        .B(shft4_w[2]), .Y(\shftOut_17[2] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_127s_8s(
       Bit_Count_16dec_i_1,
       shft2_w,
       shft1_w,
       fb_w_5,
       fb_w_0,
       fb_w_1,
       fb_w_4,
       RSControl_0_NGRST,
       N_567,
       N_570,
       N_565,
       N_569,
       N_566
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft2_w;
input  [7:0] shft1_w;
input  fb_w_5;
input  fb_w_0;
input  fb_w_1;
input  fb_w_4;
input  RSControl_0_NGRST;
input  N_567;
input  N_570;
input  N_565;
input  N_569;
input  N_566;

    wire VCC_net_1, \shftOut_8[3] , GND_net_1, \shftOut_8[4] , 
        \shftOut_8[5] , \shftOut_8[6] , \shftOut_8[7] , \shftOut_8[0] , 
        \shftOut_8[1] , \shftOut_8[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_8[5] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft2_w[5]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_8_0_a2[1]  (.A(N_567), .B(
        N_569), .C(shft1_w[1]), .D(N_566), .Y(\shftOut_8[1] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2[5]  (.A(N_570), .B(
        shft1_w[5]), .C(N_567), .Y(\shftOut_8[5] ));
    SLE \shftOut[6]  (.D(\shftOut_8[6] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft2_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_8[4] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft2_w[4]));
    SLE \shftOut[7]  (.D(\shftOut_8[7] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft2_w[7]));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2[7]  (.A(shft1_w[7]), .B(
        fb_w_5), .C(N_567), .Y(\shftOut_8[7] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_8_0_a2[0]  (.A(N_570), .B(
        shft1_w[0]), .Y(\shftOut_8[0] ));
    SLE \shftOut[3]  (.D(\shftOut_8[3] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft2_w[3]));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2[4]  (.A(N_569), .B(
        shft1_w[4]), .C(N_567), .Y(\shftOut_8[4] ));
    SLE \shftOut[2]  (.D(\shftOut_8[2] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft2_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_8[1] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft2_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_8_0_a2[3]  (.A(shft1_w[3]), .B(
        fb_w_1), .C(N_570), .Y(\shftOut_8[3] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_8_0_a2[2]  (.A(fb_w_0), .B(
        shft1_w[2]), .C(N_567), .D(N_565), .Y(\shftOut_8[2] ));
    SLE \shftOut[0]  (.D(\shftOut_8[0] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft2_w[0]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_8_0_a2[6]  (.A(fb_w_4), .B(
        shft1_w[6]), .C(N_569), .D(N_567), .Y(\shftOut_8[6] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_91s_8s(
       Bit_Count_16dec_i_1,
       shft1_w,
       shft0_w,
       fb_w_1,
       fb_w_5,
       fb_w_3,
       fb_w_0,
       fb_w_4,
       RSControl_0_NGRST,
       N_564,
       N_568,
       N_572,
       N_567,
       N_569
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft1_w;
input  [7:0] shft0_w;
input  fb_w_1;
input  fb_w_5;
input  fb_w_3;
input  fb_w_0;
input  fb_w_4;
input  RSControl_0_NGRST;
input  N_564;
input  N_568;
input  N_572;
input  N_567;
input  N_569;

    wire VCC_net_1, \shftOut_5[3] , GND_net_1, \shftOut_5[4] , 
        \shftOut_5[5] , \shftOut_5[6] , \shftOut_5[7] , \shftOut_5[0] , 
        \shftOut_5[1] , \shftOut_5[2] ;
    
    CFG2 #( .INIT(4'h6) )  \shftOut_5_0_a2[3]  (.A(N_564), .B(
        shft0_w[3]), .Y(\shftOut_5[3] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_5_0_a2[2]  (.A(fb_w_1), .B(
        shft0_w[2]), .Y(\shftOut_5[2] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_5_0_a2[6]  (.A(shft0_w[6]), .B(
        fb_w_3), .C(fb_w_5), .D(N_564), .Y(\shftOut_5[6] ));
    SLE \shftOut[5]  (.D(\shftOut_5[5] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft1_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_5[6] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft1_w[6]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \shftOut_5_0_a2[1]  (.A(shft0_w[1]), .B(
        fb_w_4), .C(fb_w_1), .D(N_569), .Y(\shftOut_5[1] ));
    SLE \shftOut[4]  (.D(\shftOut_5[4] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft1_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_5_0_a2[5]  (.A(shft0_w[5]), .B(
        fb_w_1), .C(N_572), .Y(\shftOut_5[5] ));
    SLE \shftOut[7]  (.D(\shftOut_5[7] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft1_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_5[3] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft1_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_5[2] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft1_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_5[1] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft1_w[1]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_5_0_a2[7]  (.A(shft0_w[7]), .B(
        fb_w_1), .C(fb_w_5), .D(N_572), .Y(\shftOut_5[7] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_5_0_a2[0]  (.A(shft0_w[0]), .B(
        fb_w_5), .C(N_568), .D(N_564), .Y(\shftOut_5[0] ));
    SLE \shftOut[0]  (.D(\shftOut_5[0] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft1_w[0]));
    CFG3 #( .INIT(8'h96) )  \shftOut_5_0_a2[4]  (.A(shft0_w[4]), .B(
        fb_w_0), .C(N_567), .Y(\shftOut_5[4] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_16s_8s(
       Bit_Count_16dec_i_1,
       shft4_w,
       shft3_w,
       fb_w_3,
       fb_w_4,
       fb_w_2,
       fb_w_6,
       fb_w_0,
       fb_w_7,
       fb_w_1,
       RSControl_0_NGRST,
       N_566,
       N_565
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft4_w;
input  [7:0] shft3_w;
input  fb_w_3;
input  fb_w_4;
input  fb_w_2;
input  fb_w_6;
input  fb_w_0;
input  fb_w_7;
input  fb_w_1;
input  RSControl_0_NGRST;
input  N_566;
input  N_565;

    wire VCC_net_1, \shftOut_14[3] , GND_net_1, \shftOut_14[4] , 
        \shftOut_14[5] , \shftOut_14[6] , \shftOut_14[7] , 
        \shftOut_14[0] , \shftOut_14[1] , \shftOut_14[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_14[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft4_w[5]));
    CFG2 #( .INIT(4'h6) )  \shftOut_14_0_a2[1]  (.A(fb_w_4), .B(
        shft3_w[1]), .Y(\shftOut_14[1] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_14_0_a2[0]  (.A(shft3_w[0]), .B(
        N_566), .C(N_565), .Y(\shftOut_14[0] ));
    SLE \shftOut[6]  (.D(\shftOut_14[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft4_w[6]));
    CFG3 #( .INIT(8'h96) )  \shftOut_14_0_a2[4]  (.A(fb_w_6), .B(
        shft3_w[4]), .C(fb_w_0), .Y(\shftOut_14[4] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_14[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft4_w[4]));
    CFG2 #( .INIT(4'h6) )  \shftOut_14_0_a2[3]  (.A(N_565), .B(
        shft3_w[3]), .Y(\shftOut_14[3] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_14_0_a2[2]  (.A(shft3_w[2]), .B(
        fb_w_7), .C(N_566), .Y(\shftOut_14[2] ));
    SLE \shftOut[7]  (.D(\shftOut_14[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft4_w[7]));
    CFG2 #( .INIT(4'h6) )  \shftOut_14_0_a2[6]  (.A(fb_w_2), .B(
        shft3_w[6]), .Y(\shftOut_14[6] ));
    SLE \shftOut[3]  (.D(\shftOut_14[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft4_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_14[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft4_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_14[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft4_w[1]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_14_0_a2[7]  (.A(shft3_w[7]), 
        .B(fb_w_3), .C(N_566), .D(N_565), .Y(\shftOut_14[7] ));
    SLE \shftOut[0]  (.D(\shftOut_14[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft4_w[0]));
    CFG3 #( .INIT(8'h96) )  \shftOut_14_0_a2[5]  (.A(shft3_w[5]), .B(
        fb_w_7), .C(fb_w_1), .Y(\shftOut_14[5] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_235s_8s(
       Bit_Count_16dec_i_1,
       shft7_w,
       shft6_w,
       fb_w_1,
       fb_w_6,
       fb_w_7,
       fb_w_0,
       fb_w_3,
       fb_w_5,
       fb_w_4,
       RSControl_0_NGRST,
       N_564,
       N_567
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft7_w;
input  [7:0] shft6_w;
input  fb_w_1;
input  fb_w_6;
input  fb_w_7;
input  fb_w_0;
input  fb_w_3;
input  fb_w_5;
input  fb_w_4;
input  RSControl_0_NGRST;
input  N_564;
input  N_567;

    wire VCC_net_1, \shftOut_23[3] , GND_net_1, \shftOut_23[4] , 
        \shftOut_23[5] , \shftOut_23[6] , \shftOut_23[7] , 
        \shftOut_23[0] , \shftOut_23[1] , \shftOut_23[2] ;
    
    SLE \shftOut[5]  (.D(\shftOut_23[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft7_w[5]));
    SLE \shftOut[6]  (.D(\shftOut_23[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft7_w[6]));
    CFG2 #( .INIT(4'h6) )  \shftOut_23_0_a2[5]  (.A(N_564), .B(
        shft6_w[5]), .Y(\shftOut_23[5] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_23[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft7_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_23_0_a2[3]  (.A(fb_w_7), .B(
        shft6_w[3]), .C(fb_w_0), .Y(\shftOut_23[3] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_23_0_a2[0]  (.A(shft6_w[0]), 
        .B(fb_w_4), .C(fb_w_0), .D(N_567), .Y(\shftOut_23[0] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_23_0_a2[1]  (.A(shft6_w[1]), 
        .B(fb_w_3), .C(fb_w_5), .D(N_564), .Y(\shftOut_23[1] ));
    SLE \shftOut[7]  (.D(\shftOut_23[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft7_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_23[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft7_w[3]));
    CFG2 #( .INIT(4'h6) )  \shftOut_23_0_a2[4]  (.A(fb_w_1), .B(
        shft6_w[4]), .Y(\shftOut_23[4] ));
    SLE \shftOut[2]  (.D(\shftOut_23[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft7_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_23[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft7_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_23_0_a2[6]  (.A(shft6_w[6]), .B(
        fb_w_0), .C(N_567), .Y(\shftOut_23[6] ));
    SLE \shftOut[0]  (.D(\shftOut_23[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft7_w[0]));
    CFG2 #( .INIT(4'h6) )  \shftOut_23_0_a2[2]  (.A(fb_w_6), .B(
        shft6_w[2]), .Y(\shftOut_23[2] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_23_0_a2[7]  (.A(shft6_w[7]), .B(
        fb_w_3), .C(N_564), .Y(\shftOut_23[7] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_1s_8s(
       Bit_Count_16dec_i_1,
       shft0_w,
       fb_w,
       RSControl_0_NGRST
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft0_w;
input  [7:0] fb_w;
input  RSControl_0_NGRST;

    wire VCC_net_1, GND_net_1;
    
    SLE \shftOut[4]  (.D(fb_w[4]), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft0_w[4]));
    SLE \shftOut[2]  (.D(fb_w[2]), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft0_w[2]));
    SLE \shftOut[0]  (.D(fb_w[0]), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft0_w[0]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[7]  (.D(fb_w[7]), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft0_w[7]));
    SLE \shftOut[3]  (.D(fb_w[3]), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft0_w[3]));
    SLE \shftOut[1]  (.D(fb_w[1]), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft0_w[1]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[5]  (.D(fb_w[5]), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft0_w[5]));
    SLE \shftOut[6]  (.D(fb_w[6]), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(shft0_w[6]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_54s_8s_0(
       Bit_Count_16dec_i_1,
       shft20_w,
       shft19_w,
       fb_w_3,
       fb_w_0,
       fb_w_5,
       fb_w_2,
       fb_w_1,
       fb_w_7,
       RSControl_0_NGRST,
       N_588,
       N_568,
       N_575,
       N_566,
       N_573,
       N_567,
       N_569,
       N_572,
       N_565
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft20_w;
input  [7:0] shft19_w;
input  fb_w_3;
input  fb_w_0;
input  fb_w_5;
input  fb_w_2;
input  fb_w_1;
input  fb_w_7;
input  RSControl_0_NGRST;
output N_588;
input  N_568;
input  N_575;
input  N_566;
input  N_573;
input  N_567;
input  N_569;
input  N_572;
input  N_565;

    wire VCC_net_1, \shftOut_38[3] , GND_net_1, \shftOut_38[4] , 
        \shftOut_38[5] , \shftOut_38[6] , \shftOut_38[7] , 
        \shftOut_38[0] , \shftOut_38[1] , \shftOut_38[2] ;
    
    CFG2 #( .INIT(4'h6) )  \shftOut_38_0_a2_0[1]  (.A(fb_w_3), .B(
        fb_w_0), .Y(N_588));
    SLE \shftOut[5]  (.D(\shftOut_38[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft20_w[5]));
    CFG3 #( .INIT(8'h96) )  \shftOut_38_0_a2[7]  (.A(fb_w_5), .B(
        shft19_w[7]), .C(fb_w_2), .Y(\shftOut_38[7] ));
    SLE \shftOut[6]  (.D(\shftOut_38[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft20_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_38[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft20_w[4]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_38_0_a2[5]  (.A(shft19_w[5]), 
        .B(fb_w_0), .C(N_575), .D(N_566), .Y(\shftOut_38[5] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_38_0_a2[4]  (.A(N_569), .B(
        shft19_w[4]), .C(N_568), .Y(\shftOut_38[4] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_38_0_a2[3]  (.A(shft19_w[3]), 
        .B(fb_w_2), .C(fb_w_1), .D(N_573), .Y(\shftOut_38[3] ));
    SLE \shftOut[7]  (.D(\shftOut_38[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft20_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_38[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft20_w[3]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_38_0_a2[6]  (.A(shft19_w[6]), 
        .B(fb_w_1), .C(N_572), .D(N_565), .Y(\shftOut_38[6] ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_38_0_a2[2]  (.A(fb_w_0), .B(
        shft19_w[2]), .C(N_573), .D(N_567), .Y(\shftOut_38[2] ));
    SLE \shftOut[2]  (.D(\shftOut_38[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft20_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_38[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft20_w[1]));
    CFG2 #( .INIT(4'h6) )  \shftOut_38_0_a2[0]  (.A(N_568), .B(
        shft19_w[0]), .Y(\shftOut_38[0] ));
    SLE \shftOut[0]  (.D(\shftOut_38[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft20_w[0]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_38_0_a2[1]  (.A(shft19_w[1]), 
        .B(fb_w_7), .C(N_588), .D(N_566), .Y(\shftOut_38[1] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_8s_8s(
       Bit_Count_16dec_i_1,
       shft10_w,
       shft9_w,
       fb_w_2,
       fb_w_5,
       fb_w_3,
       fb_w_6,
       fb_w_0,
       fb_w_7,
       fb_w_1,
       RSControl_0_NGRST,
       N_566,
       N_565
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft10_w;
input  [7:0] shft9_w;
input  fb_w_2;
input  fb_w_5;
input  fb_w_3;
input  fb_w_6;
input  fb_w_0;
input  fb_w_7;
input  fb_w_1;
input  RSControl_0_NGRST;
input  N_566;
input  N_565;

    wire VCC_net_1, \shftOut_32[3] , GND_net_1, \shftOut_32[4] , 
        \shftOut_32[5] , \shftOut_32[6] , \shftOut_32[7] , 
        \shftOut_32[0] , \shftOut_32[1] , \shftOut_32[2] ;
    
    CFG3 #( .INIT(8'h96) )  \shftOut_32_0_a2[0]  (.A(shft9_w[0]), .B(
        fb_w_6), .C(N_565), .Y(\shftOut_32[0] ));
    SLE \shftOut[5]  (.D(\shftOut_32[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft10_w[5]));
    CFG2 #( .INIT(4'h6) )  \shftOut_32_0_a2[1]  (.A(fb_w_5), .B(
        shft9_w[1]), .Y(\shftOut_32[1] ));
    SLE \shftOut[6]  (.D(\shftOut_32[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft10_w[6]));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_32[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft10_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_32_0_a2[7]  (.A(shft9_w[7]), .B(
        N_566), .C(N_565), .Y(\shftOut_32[7] ));
    SLE \shftOut[7]  (.D(\shftOut_32[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft10_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_32[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft10_w[3]));
    CFG2 #( .INIT(4'h6) )  \shftOut_32_0_a2[5]  (.A(fb_w_2), .B(
        shft9_w[5]), .Y(\shftOut_32[5] ));
    SLE \shftOut[2]  (.D(\shftOut_32[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft10_w[2]));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'h96) )  \shftOut_32_0_a2[4]  (.A(shft9_w[4]), .B(
        fb_w_7), .C(fb_w_1), .Y(\shftOut_32[4] ));
    SLE \shftOut[1]  (.D(\shftOut_32[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft10_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_32_0_a2[3]  (.A(fb_w_6), .B(
        shft9_w[3]), .C(fb_w_0), .Y(\shftOut_32[3] ));
    SLE \shftOut[0]  (.D(\shftOut_32[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft10_w[0]));
    CFG2 #( .INIT(4'h6) )  \shftOut_32_0_a2[6]  (.A(fb_w_3), .B(
        shft9_w[6]), .Y(\shftOut_32[6] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_32_0_a2[2]  (.A(N_565), .B(
        shft9_w[2]), .Y(\shftOut_32[2] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_lastTap_91s_8s(
       Bit_Count_16dec_i_1,
       dInp_reg_w,
       parity_w,
       pre_fb_w,
       conv_basis,
       fb_w,
       shft30_w,
       RSControl_0_NGRST,
       hold0fb_w,
       N_564,
       N_569,
       N_572,
       N_568,
       N_567
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] dInp_reg_w;
output [7:0] parity_w;
output [7:0] pre_fb_w;
input  [7:0] conv_basis;
input  [7:0] fb_w;
input  [7:0] shft30_w;
input  RSControl_0_NGRST;
input  hold0fb_w;
output N_564;
output N_569;
output N_572;
output N_568;
input  N_567;

    wire VCC_net_1, \shftOut_2[2] , GND_net_1, \shftOut_2[3] , 
        \shftOut_2[4] , \shftOut_2[5] , \shftOut_2[6] , \shftOut_2[7] , 
        \pre_fbOut_4[3]_net_1 , \pre_fbOut_4[4]_net_1 , 
        \pre_fbOut_4[5]_net_1 , \pre_fbOut_4[6]_net_1 , 
        \pre_fbOut_4[7]_net_1 , \dInp_reg_4[0]_net_1 , 
        \dInp_reg_4[1]_net_1 , \dInp_reg_4[2]_net_1 , 
        \dInp_reg_4[3]_net_1 , \dInp_reg_4[4]_net_1 , 
        \dInp_reg_4[5]_net_1 , \dInp_reg_4[6]_net_1 , 
        \dInp_reg_4[7]_net_1 , \shftOut_2[0] , \shftOut_2[1] , 
        \pre_fbOut_4[0]_net_1 , \pre_fbOut_4[1]_net_1 , 
        \pre_fbOut_4[2]_net_1 ;
    
    SLE \pre_fbOut[2]  (.D(\pre_fbOut_4[2]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(pre_fb_w[2]));
    CFG2 #( .INIT(4'h4) )  \dInp_reg_4[6]  (.A(hold0fb_w), .B(
        conv_basis[6]), .Y(\dInp_reg_4[6]_net_1 ));
    SLE \shftOut[3]  (.D(\shftOut_2[3] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(parity_w[3]));
    SLE \dInp_reg[4]  (.D(\dInp_reg_4[4]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dInp_reg_w[4]));
    CFG2 #( .INIT(4'h2) )  \pre_fbOut_4[2]  (.A(\shftOut_2[2] ), .B(
        hold0fb_w), .Y(\pre_fbOut_4[2]_net_1 ));
    SLE \shftOut[0]  (.D(\shftOut_2[0] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(parity_w[0]));
    SLE \pre_fbOut[7]  (.D(\pre_fbOut_4[7]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(pre_fb_w[7]));
    SLE \shftOut[2]  (.D(\shftOut_2[2] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(parity_w[2]));
    SLE \dInp_reg[3]  (.D(\dInp_reg_4[3]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dInp_reg_w[3]));
    CFG2 #( .INIT(4'h2) )  \pre_fbOut_4[7]  (.A(\shftOut_2[7] ), .B(
        hold0fb_w), .Y(\pre_fbOut_4[7]_net_1 ));
    SLE \pre_fbOut[1]  (.D(\pre_fbOut_4[1]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(pre_fb_w[1]));
    CFG3 #( .INIT(8'h96) )  \shftOut_2_0_a2[5]  (.A(shft30_w[5]), .B(
        fb_w[1]), .C(N_572), .Y(\shftOut_2[5] ));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[6]  (.D(\shftOut_2[6] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(parity_w[6]));
    SLE \pre_fbOut[5]  (.D(\pre_fbOut_4[5]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(pre_fb_w[5]));
    CFG2 #( .INIT(4'h2) )  \pre_fbOut_4[1]  (.A(\shftOut_2[1] ), .B(
        hold0fb_w), .Y(\pre_fbOut_4[1]_net_1 ));
    SLE \shftOut[7]  (.D(\shftOut_2[7] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(parity_w[7]));
    SLE \shftOut[5]  (.D(\shftOut_2[5] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(parity_w[5]));
    CFG3 #( .INIT(8'h14) )  \pre_fbOut_4[3]  (.A(hold0fb_w), .B(N_564), 
        .C(shft30_w[3]), .Y(\pre_fbOut_4[3]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_2_0_a2[0]  (.A(shft30_w[0]), 
        .B(fb_w[5]), .C(N_568), .D(N_564), .Y(\shftOut_2[0] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_2_0_a2_0[0]  (.A(fb_w[3]), .B(
        fb_w[6]), .Y(N_568));
    SLE \pre_fbOut[3]  (.D(\pre_fbOut_4[3]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(pre_fb_w[3]));
    CFG2 #( .INIT(4'h4) )  \dInp_reg_4[4]  (.A(hold0fb_w), .B(
        conv_basis[4]), .Y(\dInp_reg_4[4]_net_1 ));
    SLE \dInp_reg[2]  (.D(\dInp_reg_4[2]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dInp_reg_w[2]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \shftOut_2_0_a2[1]  (.A(shft30_w[1]), 
        .B(fb_w[4]), .C(fb_w[1]), .D(N_569), .Y(\shftOut_2[1] ));
    CFG2 #( .INIT(4'h4) )  \dInp_reg_4[2]  (.A(hold0fb_w), .B(
        conv_basis[2]), .Y(\dInp_reg_4[2]_net_1 ));
    SLE \shftOut[4]  (.D(\shftOut_2[4] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(parity_w[4]));
    SLE \dInp_reg[6]  (.D(\dInp_reg_4[6]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dInp_reg_w[6]));
    CFG2 #( .INIT(4'h6) )  \shftOut_2_0_a2[2]  (.A(fb_w[1]), .B(
        shft30_w[2]), .Y(\shftOut_2[2] ));
    SLE \pre_fbOut[4]  (.D(\pre_fbOut_4[4]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(pre_fb_w[4]));
    SLE \dInp_reg[7]  (.D(\dInp_reg_4[7]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dInp_reg_w[7]));
    CFG2 #( .INIT(4'h2) )  \pre_fbOut_4[4]  (.A(\shftOut_2[4] ), .B(
        hold0fb_w), .Y(\pre_fbOut_4[4]_net_1 ));
    SLE \dInp_reg[1]  (.D(\dInp_reg_4[1]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dInp_reg_w[1]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_2_0_a2[7]  (.A(shft30_w[7]), 
        .B(fb_w[1]), .C(fb_w[5]), .D(N_572), .Y(\shftOut_2[7] ));
    SLE \pre_fbOut[6]  (.D(\pre_fbOut_4[6]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(pre_fb_w[6]));
    SLE \shftOut[1]  (.D(\shftOut_2[1] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(parity_w[1]));
    CFG2 #( .INIT(4'h2) )  \pre_fbOut_4[6]  (.A(\shftOut_2[6] ), .B(
        hold0fb_w), .Y(\pre_fbOut_4[6]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \shftOut_2_0_a2[3]  (.A(N_564), .B(
        shft30_w[3]), .Y(\shftOut_2[3] ));
    SLE \dInp_reg[5]  (.D(\dInp_reg_4[5]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dInp_reg_w[5]));
    CFG3 #( .INIT(8'h96) )  \shftOut_2_0_a2_0[3]  (.A(dInp_reg_w[2]), 
        .B(fb_w[0]), .C(pre_fb_w[2]), .Y(N_564));
    CFG2 #( .INIT(4'h4) )  \dInp_reg_4[5]  (.A(hold0fb_w), .B(
        conv_basis[5]), .Y(\dInp_reg_4[5]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \pre_fbOut_4[5]  (.A(\shftOut_2[5] ), .B(
        hold0fb_w), .Y(\pre_fbOut_4[5]_net_1 ));
    SLE \pre_fbOut[0]  (.D(\pre_fbOut_4[0]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(pre_fb_w[0]));
    CFG2 #( .INIT(4'h4) )  \dInp_reg_4[7]  (.A(hold0fb_w), .B(
        conv_basis[7]), .Y(\dInp_reg_4[7]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \dInp_reg_4[0]  (.A(hold0fb_w), .B(
        conv_basis[0]), .Y(\dInp_reg_4[0]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  \shftOut_2_0_a2_0[1]  (.A(fb_w[7]), .B(
        N_564), .C(pre_fb_w[5]), .D(dInp_reg_w[5]), .Y(N_569));
    CFG2 #( .INIT(4'h2) )  \pre_fbOut_4[0]  (.A(\shftOut_2[0] ), .B(
        hold0fb_w), .Y(\pre_fbOut_4[0]_net_1 ));
    CFG3 #( .INIT(8'h96) )  \shftOut_2_0_a2[4]  (.A(shft30_w[4]), .B(
        fb_w[0]), .C(N_567), .Y(\shftOut_2[4] ));
    CFG2 #( .INIT(4'h4) )  \dInp_reg_4[3]  (.A(hold0fb_w), .B(
        conv_basis[3]), .Y(\dInp_reg_4[3]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \shftOut_2_0_a2_0[7]  (.A(fb_w[2]), .B(
        fb_w[4]), .Y(N_572));
    CFG4 #( .INIT(16'h6996) )  \shftOut_2_0_a2[6]  (.A(shft30_w[6]), 
        .B(fb_w[3]), .C(fb_w[5]), .D(N_564), .Y(\shftOut_2[6] ));
    CFG2 #( .INIT(4'h4) )  \dInp_reg_4[1]  (.A(hold0fb_w), .B(
        conv_basis[1]), .Y(\dInp_reg_4[1]_net_1 ));
    SLE \dInp_reg[0]  (.D(\dInp_reg_4[0]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(dInp_reg_w[0]));
    
endmodule


module TM_RSENC_TM_RSENC_0_rsEnc_tap_13s_8s(
       Bit_Count_16dec_i_1,
       shft6_w,
       shft5_w,
       fb_w_5,
       fb_w_3,
       fb_w_2,
       fb_w_7,
       fb_w_1,
       fb_w_0,
       fb_w_6,
       RSControl_0_NGRST,
       N_576,
       N_583,
       N_574,
       N_566,
       N_572,
       N_575,
       N_569
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] shft6_w;
input  [7:0] shft5_w;
input  fb_w_5;
input  fb_w_3;
input  fb_w_2;
input  fb_w_7;
input  fb_w_1;
input  fb_w_0;
input  fb_w_6;
input  RSControl_0_NGRST;
input  N_576;
input  N_583;
input  N_574;
input  N_566;
input  N_572;
input  N_575;
input  N_569;

    wire VCC_net_1, \shftOut_20[3] , GND_net_1, \shftOut_20[4] , 
        \shftOut_20[5] , \shftOut_20[6] , \shftOut_20[7] , 
        \shftOut_20[0] , \shftOut_20[1] , \shftOut_20[2] ;
    
    CFG2 #( .INIT(4'h6) )  \shftOut_20_0_a2[0]  (.A(N_583), .B(
        shft5_w[0]), .Y(\shftOut_20[0] ));
    SLE \shftOut[5]  (.D(\shftOut_20[5] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft6_w[5]));
    CFG3 #( .INIT(8'h96) )  \shftOut_20_0_a2[1]  (.A(shft5_w[1]), .B(
        fb_w_5), .C(N_574), .Y(\shftOut_20[1] ));
    SLE \shftOut[6]  (.D(\shftOut_20[6] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft6_w[6]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_20_0_a2[4]  (.A(shft5_w[4]), 
        .B(fb_w_7), .C(fb_w_1), .D(N_572), .Y(\shftOut_20[4] ));
    GND GND (.Y(GND_net_1));
    SLE \shftOut[4]  (.D(\shftOut_20[4] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft6_w[4]));
    CFG3 #( .INIT(8'h96) )  \shftOut_20_0_a2[6]  (.A(shft5_w[6]), .B(
        fb_w_3), .C(N_566), .Y(\shftOut_20[6] ));
    CFG3 #( .INIT(8'h96) )  \shftOut_20_0_a2[2]  (.A(shft5_w[2]), .B(
        fb_w_6), .C(N_569), .Y(\shftOut_20[2] ));
    CFG2 #( .INIT(4'h6) )  \shftOut_20_0_a2[7]  (.A(N_576), .B(
        shft5_w[7]), .Y(\shftOut_20[7] ));
    SLE \shftOut[7]  (.D(\shftOut_20[7] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft6_w[7]));
    SLE \shftOut[3]  (.D(\shftOut_20[3] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft6_w[3]));
    SLE \shftOut[2]  (.D(\shftOut_20[2] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft6_w[2]));
    VCC VCC (.Y(VCC_net_1));
    SLE \shftOut[1]  (.D(\shftOut_20[1] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft6_w[1]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_20_0_a2[5]  (.A(fb_w_3), .B(
        fb_w_5), .C(shft5_w[5]), .D(fb_w_2), .Y(\shftOut_20[5] ));
    SLE \shftOut[0]  (.D(\shftOut_20[0] ), .CLK(Bit_Count_16dec_i_1[3])
        , .EN(VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shft6_w[0]));
    CFG4 #( .INIT(16'h6996) )  \shftOut_20_0_a2[3]  (.A(shft5_w[3]), 
        .B(fb_w_0), .C(fb_w_6), .D(N_575), .Y(\shftOut_20[3] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_gfIIR_8s(
       Bit_Count_16dec_i_1,
       encoded,
       conv_basis,
       RSControl_0_NGRST,
       datNotParity_w,
       hold0fb_w
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] encoded;
input  [7:0] conv_basis;
input  RSControl_0_NGRST;
input  datNotParity_w;
input  hold0fb_w;

    wire VCC_net_1, \codeOut_3[0]_net_1 , GND_net_1, 
        \codeOut_3[1]_net_1 , \codeOut_3[2]_net_1 , 
        \codeOut_3[3]_net_1 , \codeOut_3[4]_net_1 , 
        \codeOut_3[5]_net_1 , \codeOut_3[6]_net_1 , 
        \codeOut_3[7]_net_1 , \dInp_reg_w[1] , \pre_fb_w[1] , 
        \fb_w[1] , \dInp_reg_w[7] , \pre_fb_w[7] , \fb_w[7] , 
        \dInp_reg_w[0] , \pre_fb_w[0] , \fb_w[0] , \dInp_reg_w[4] , 
        \pre_fb_w[4] , \fb_w[4] , \dInp_reg_w[2] , \pre_fb_w[2] , 
        \fb_w[2] , \dInp_reg_w[5] , \pre_fb_w[5] , \fb_w[5] , 
        \dInp_reg_w[3] , \pre_fb_w[3] , \fb_w[3] , \dInp_reg_w[6] , 
        \pre_fb_w[6] , \fb_w[6] , \parity_w[0] , \parity_w[1] , 
        \parity_w[2] , \parity_w[3] , \parity_w[5] , \parity_w[7] , 
        \parity_w[6] , \parity_w[4] , \shft0_w[0] , \shft0_w[1] , 
        \shft0_w[2] , \shft0_w[3] , \shft0_w[4] , \shft0_w[5] , 
        \shft0_w[6] , \shft0_w[7] , \shft1_w[0] , \shft1_w[1] , 
        \shft1_w[2] , \shft1_w[3] , \shft1_w[4] , \shft1_w[5] , 
        \shft1_w[6] , \shft1_w[7] , N_564, N_568, N_572, N_567, N_569, 
        \shft2_w[0] , \shft2_w[1] , \shft2_w[2] , \shft2_w[3] , 
        \shft2_w[4] , \shft2_w[5] , \shft2_w[6] , \shft2_w[7] , N_570, 
        N_565, N_566, \shft3_w[0] , \shft3_w[1] , \shft3_w[2] , 
        \shft3_w[3] , \shft3_w[4] , \shft3_w[5] , \shft3_w[6] , 
        \shft3_w[7] , N_574, N_576, N_575, \shft4_w[0] , \shft4_w[1] , 
        \shft4_w[2] , \shft4_w[3] , \shft4_w[4] , \shft4_w[5] , 
        \shft4_w[6] , \shft4_w[7] , \shft5_w[0] , \shft5_w[1] , 
        \shft5_w[2] , \shft5_w[3] , \shft5_w[4] , \shft5_w[5] , 
        \shft5_w[6] , \shft5_w[7] , \shftOut_17_1[2] , \shft6_w[0] , 
        \shft6_w[1] , \shft6_w[2] , \shft6_w[3] , \shft6_w[4] , 
        \shft6_w[5] , \shft6_w[6] , \shft6_w[7] , N_583, \shft7_w[0] , 
        \shft7_w[1] , \shft7_w[2] , \shft7_w[3] , \shft7_w[4] , 
        \shft7_w[5] , \shft7_w[6] , \shft7_w[7] , \shft8_w[0] , 
        \shft8_w[1] , \shft8_w[2] , \shft8_w[3] , \shft8_w[4] , 
        \shft8_w[5] , \shft8_w[6] , \shft8_w[7] , \shft9_w[0] , 
        \shft9_w[1] , \shft9_w[2] , \shft9_w[3] , \shft9_w[4] , 
        \shft9_w[5] , \shft9_w[6] , \shft9_w[7] , N_588, \shft10_w[0] , 
        \shft10_w[1] , \shft10_w[2] , \shft10_w[3] , \shft10_w[4] , 
        \shft10_w[5] , \shft10_w[6] , \shft10_w[7] , \shft11_w[0] , 
        \shft11_w[1] , \shft11_w[2] , \shft11_w[3] , \shft11_w[4] , 
        \shft11_w[5] , \shft11_w[6] , \shft11_w[7] , \shft12_w[0] , 
        \shft12_w[1] , \shft12_w[2] , \shft12_w[3] , \shft12_w[4] , 
        \shft12_w[5] , \shft12_w[6] , \shft12_w[7] , N_573, 
        \shft13_w[0] , \shft13_w[1] , \shft13_w[2] , \shft13_w[3] , 
        \shft13_w[4] , \shft13_w[5] , \shft13_w[6] , \shft13_w[7] , 
        \shft14_w[0] , \shft14_w[1] , \shft14_w[2] , \shft14_w[3] , 
        \shft14_w[4] , \shft14_w[5] , \shft14_w[6] , \shft14_w[7] , 
        \shft15_w[0] , \shft15_w[1] , \shft15_w[2] , \shft15_w[3] , 
        \shft15_w[4] , \shft15_w[5] , \shft15_w[6] , \shft15_w[7] , 
        \shft16_w[0] , \shft16_w[1] , \shft16_w[2] , \shft16_w[3] , 
        \shft16_w[4] , \shft16_w[5] , \shft16_w[6] , \shft16_w[7] , 
        \shft17_w[0] , \shft17_w[1] , \shft17_w[2] , \shft17_w[3] , 
        \shft17_w[4] , \shft17_w[5] , \shft17_w[6] , \shft17_w[7] , 
        \shft18_w[0] , \shft18_w[1] , \shft18_w[2] , \shft18_w[3] , 
        \shft18_w[4] , \shft18_w[5] , \shft18_w[6] , \shft18_w[7] , 
        \shft19_w[0] , \shft19_w[1] , \shft19_w[2] , \shft19_w[3] , 
        \shft19_w[4] , \shft19_w[5] , \shft19_w[6] , \shft19_w[7] , 
        \shft20_w[0] , \shft20_w[1] , \shft20_w[2] , \shft20_w[3] , 
        \shft20_w[4] , \shft20_w[5] , \shft20_w[6] , \shft20_w[7] , 
        \shft21_w[0] , \shft21_w[1] , \shft21_w[2] , \shft21_w[3] , 
        \shft21_w[4] , \shft21_w[5] , \shft21_w[6] , \shft21_w[7] , 
        \shft22_w[0] , \shft22_w[1] , \shft22_w[2] , \shft22_w[3] , 
        \shft22_w[4] , \shft22_w[5] , \shft22_w[6] , \shft22_w[7] , 
        \shft23_w[0] , \shft23_w[1] , \shft23_w[2] , \shft23_w[3] , 
        \shft23_w[4] , \shft23_w[5] , \shft23_w[6] , \shft23_w[7] , 
        \shft24_w[0] , \shft24_w[1] , \shft24_w[2] , \shft24_w[3] , 
        \shft24_w[4] , \shft24_w[5] , \shft24_w[6] , \shft24_w[7] , 
        \shft25_w[0] , \shft25_w[1] , \shft25_w[2] , \shft25_w[3] , 
        \shft25_w[4] , \shft25_w[5] , \shft25_w[6] , \shft25_w[7] , 
        \shft26_w[0] , \shft26_w[1] , \shft26_w[2] , \shft26_w[3] , 
        \shft26_w[4] , \shft26_w[5] , \shft26_w[6] , \shft26_w[7] , 
        \shft27_w[0] , \shft27_w[1] , \shft27_w[2] , \shft27_w[3] , 
        \shft27_w[4] , \shft27_w[5] , \shft27_w[6] , \shft27_w[7] , 
        \shft28_w[0] , \shft28_w[1] , \shft28_w[2] , \shft28_w[3] , 
        \shft28_w[4] , \shft28_w[5] , \shft28_w[6] , \shft28_w[7] , 
        \shft29_w[0] , \shft29_w[1] , \shft29_w[2] , \shft29_w[3] , 
        \shft29_w[4] , \shft29_w[5] , \shft29_w[6] , \shft29_w[7] , 
        \shft30_w[0] , \shft30_w[1] , \shft30_w[2] , \shft30_w[3] , 
        \shft30_w[4] , \shft30_w[5] , \shft30_w[6] , \shft30_w[7] ;
    
    CFG3 #( .INIT(8'hCA) )  \codeOut_3[7]  (.A(\parity_w[7] ), .B(
        \dInp_reg_w[7] ), .C(datNotParity_w), .Y(\codeOut_3[7]_net_1 ));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_165s_8s tap_9 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft9_w({\shft9_w[7] , \shft9_w[6] , 
        \shft9_w[5] , \shft9_w[4] , \shft9_w[3] , \shft9_w[2] , 
        \shft9_w[1] , \shft9_w[0] }), .shft8_w({\shft8_w[7] , 
        \shft8_w[6] , \shft8_w[5] , \shft8_w[4] , \shft8_w[3] , 
        \shft8_w[2] , \shft8_w[1] , \shft8_w[0] }), .fb_w_1(\fb_w[1] ), 
        .fb_w_5(\fb_w[5] ), .fb_w_7(\fb_w[7] ), .fb_w_2(\fb_w[2] ), 
        .fb_w_0(\fb_w[0] ), .fb_w_4(\fb_w[4] ), .fb_w_3(\fb_w[3] ), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_566(N_566), .N_568(
        N_568), .N_574(N_574), .N_564(N_564), .N_570(N_570), .N_567(
        N_567), .N_565(N_565), .N_588(N_588));
    CFG3 #( .INIT(8'hCA) )  \codeOut_3[3]  (.A(\parity_w[3] ), .B(
        \dInp_reg_w[3] ), .C(datNotParity_w), .Y(\codeOut_3[3]_net_1 ));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_86s_8s_2 tap_29 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft29_w({
        \shft29_w[7] , \shft29_w[6] , \shft29_w[5] , \shft29_w[4] , 
        \shft29_w[3] , \shft29_w[2] , \shft29_w[1] , \shft29_w[0] }), 
        .shft28_w({\shft28_w[7] , \shft28_w[6] , \shft28_w[5] , 
        \shft28_w[4] , \shft28_w[3] , \shft28_w[2] , \shft28_w[1] , 
        \shft28_w[0] }), .fb_w({\fb_w[7] , \fb_w[6] , \fb_w[5] , 
        \fb_w[4] , \fb_w[3] , \fb_w[2] , \fb_w[1] }), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_568(N_568), .N_567(
        N_567), .N_574(N_574), .N_569(N_569), .N_576(N_576), .N_564(
        N_564), .N_565(N_565), .N_570(N_570), .N_575(N_575));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_86s_8s_1 tap_19 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft19_w({
        \shft19_w[7] , \shft19_w[6] , \shft19_w[5] , \shft19_w[4] , 
        \shft19_w[3] , \shft19_w[2] , \shft19_w[1] , \shft19_w[0] }), 
        .shft18_w({\shft18_w[7] , \shft18_w[6] , \shft18_w[5] , 
        \shft18_w[4] , \shft18_w[3] , \shft18_w[2] , \shft18_w[1] , 
        \shft18_w[0] }), .fb_w({\fb_w[7] , \fb_w[6] , \fb_w[5] , 
        \fb_w[4] , \fb_w[3] , \fb_w[2] , \fb_w[1] }), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_568(N_568), .N_567(
        N_567), .N_574(N_574), .N_569(N_569), .N_576(N_576), .N_564(
        N_564), .N_565(N_565), .N_570(N_570), .N_575(N_575));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_86s_8s tap_3 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft3_w({\shft3_w[7] , \shft3_w[6] , 
        \shft3_w[5] , \shft3_w[4] , \shft3_w[3] , \shft3_w[2] , 
        \shft3_w[1] , \shft3_w[0] }), .shft2_w({\shft2_w[7] , 
        \shft2_w[6] , \shft2_w[5] , \shft2_w[4] , \shft2_w[3] , 
        \shft2_w[2] , \shft2_w[1] , \shft2_w[0] }), .fb_w({\fb_w[7] , 
        \fb_w[6] , \fb_w[5] , \fb_w[4] , \fb_w[3] , \fb_w[2] , 
        \fb_w[1] }), .RSControl_0_NGRST(RSControl_0_NGRST), .N_568(
        N_568), .N_567(N_567), .N_574(N_574), .N_569(N_569), .N_576(
        N_576), .N_564(N_564), .N_565(N_565), .N_570(N_570), .N_575(
        N_575));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_30s_8s_0 tap_27 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft27_w({
        \shft27_w[7] , \shft27_w[6] , \shft27_w[5] , \shft27_w[4] , 
        \shft27_w[3] , \shft27_w[2] , \shft27_w[1] , \shft27_w[0] }), 
        .pre_fb_w({\pre_fb_w[3] }), .dInp_reg_w({\dInp_reg_w[3] }), 
        .shftOut_17_1({\shftOut_17_1[2] }), .shft26_w({\shft26_w[7] , 
        \shft26_w[6] , \shft26_w[5] , \shft26_w[4] , \shft26_w[3] , 
        \shft26_w[2] , \shft26_w[1] , \shft26_w[0] }), .fb_w_0(
        \fb_w[0] ), .fb_w_7(\fb_w[7] ), .fb_w_1(\fb_w[1] ), .fb_w_5(
        \fb_w[5] ), .fb_w_3(\fb_w[3] ), .fb_w_4(\fb_w[4] ), .fb_w_6(
        \fb_w[6] ), .RSControl_0_NGRST(RSControl_0_NGRST), .N_566(
        N_566), .N_565(N_565), .N_575(N_575), .N_572(N_572), .N_574(
        N_574), .N_564(N_564));
    CFG2 #( .INIT(4'h6) )  \fb_w_i_o2[3]  (.A(\dInp_reg_w[3] ), .B(
        \pre_fb_w[3] ), .Y(\fb_w[3] ));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_32s_8s_0 tap_17 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft17_w({
        \shft17_w[7] , \shft17_w[6] , \shft17_w[5] , \shft17_w[4] , 
        \shft17_w[3] , \shft17_w[2] , \shft17_w[1] , \shft17_w[0] }), 
        .shft16_w({\shft16_w[7] , \shft16_w[6] , \shft16_w[5] , 
        \shft16_w[4] , \shft16_w[3] , \shft16_w[2] , \shft16_w[1] , 
        \shft16_w[0] }), .fb_w_3(\fb_w[3] ), .fb_w_6(\fb_w[6] ), 
        .fb_w_0(\fb_w[0] ), .fb_w_7(\fb_w[7] ), .fb_w_1(\fb_w[1] ), 
        .fb_w_2(\fb_w[2] ), .RSControl_0_NGRST(RSControl_0_NGRST), 
        .N_566(N_566), .N_565(N_565), .N_568(N_568), .N_573(N_573));
    CFG3 #( .INIT(8'hCA) )  \codeOut_3[6]  (.A(\parity_w[6] ), .B(
        \dInp_reg_w[6] ), .C(datNotParity_w), .Y(\codeOut_3[6]_net_1 ));
    SLE \codeOut[2]  (.D(\codeOut_3[2]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(encoded[2]));
    SLE \codeOut[4]  (.D(\codeOut_3[4]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(encoded[4]));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_16s_8s_0 tap_28 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft28_w({
        \shft28_w[7] , \shft28_w[6] , \shft28_w[5] , \shft28_w[4] , 
        \shft28_w[3] , \shft28_w[2] , \shft28_w[1] , \shft28_w[0] }), 
        .shft27_w({\shft27_w[7] , \shft27_w[6] , \shft27_w[5] , 
        \shft27_w[4] , \shft27_w[3] , \shft27_w[2] , \shft27_w[1] , 
        \shft27_w[0] }), .fb_w_3(\fb_w[3] ), .fb_w_4(\fb_w[4] ), 
        .fb_w_2(\fb_w[2] ), .fb_w_6(\fb_w[6] ), .fb_w_0(\fb_w[0] ), 
        .fb_w_7(\fb_w[7] ), .fb_w_1(\fb_w[1] ), .RSControl_0_NGRST(
        RSControl_0_NGRST), .N_566(N_566), .N_565(N_565), .N_573(N_573)
        );
    TM_RSENC_TM_RSENC_0_rsEnc_tap_171s_8s_0 tap_18 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft18_w({
        \shft18_w[7] , \shft18_w[6] , \shft18_w[5] , \shft18_w[4] , 
        \shft18_w[3] , \shft18_w[2] , \shft18_w[1] , \shft18_w[0] }), 
        .shft17_w({\shft17_w[7] , \shft17_w[6] , \shft17_w[5] , 
        \shft17_w[4] , \shft17_w[3] , \shft17_w[2] , \shft17_w[1] , 
        \shft17_w[0] }), .fb_w_1(\fb_w[1] ), .fb_w_7(\fb_w[7] ), 
        .fb_w_3(\fb_w[3] ), .fb_w_5(\fb_w[5] ), .fb_w_0(\fb_w[0] ), 
        .fb_w_6(\fb_w[6] ), .RSControl_0_NGRST(RSControl_0_NGRST), 
        .N_583(N_583), .N_566(N_566), .N_569(N_569), .N_568(N_568), 
        .N_572(N_572), .N_565(N_565), .N_567(N_567), .N_574(N_574));
    SLE \codeOut[7]  (.D(\codeOut_3[7]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(encoded[7]));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_97s_8s tap_8 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft8_w({\shft8_w[7] , \shft8_w[6] , 
        \shft8_w[5] , \shft8_w[4] , \shft8_w[3] , \shft8_w[2] , 
        \shft8_w[1] , \shft8_w[0] }), .shft7_w({\shft7_w[7] , 
        \shft7_w[6] , \shft7_w[5] , \shft7_w[4] , \shft7_w[3] , 
        \shft7_w[2] , \shft7_w[1] , \shft7_w[0] }), .fb_w({\fb_w[7] , 
        \fb_w[6] , \fb_w[5] , \fb_w[4] , \fb_w[3] , \fb_w[2] , 
        \fb_w[1] , \fb_w[0] }), .RSControl_0_NGRST(RSControl_0_NGRST), 
        .N_564(N_564), .N_567(N_567));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_235s_8s_0 tap_25 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft25_w({
        \shft25_w[7] , \shft25_w[6] , \shft25_w[5] , \shft25_w[4] , 
        \shft25_w[3] , \shft25_w[2] , \shft25_w[1] , \shft25_w[0] }), 
        .shft24_w({\shft24_w[7] , \shft24_w[6] , \shft24_w[5] , 
        \shft24_w[4] , \shft24_w[3] , \shft24_w[2] , \shft24_w[1] , 
        \shft24_w[0] }), .fb_w_1(\fb_w[1] ), .fb_w_6(\fb_w[6] ), 
        .fb_w_7(\fb_w[7] ), .fb_w_0(\fb_w[0] ), .fb_w_3(\fb_w[3] ), 
        .fb_w_5(\fb_w[5] ), .fb_w_4(\fb_w[4] ), .RSControl_0_NGRST(
        RSControl_0_NGRST), .N_564(N_564), .N_567(N_567));
    VCC VCC (.Y(VCC_net_1));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_32s_8s tap_15 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft15_w({\shft15_w[7] , 
        \shft15_w[6] , \shft15_w[5] , \shft15_w[4] , \shft15_w[3] , 
        \shft15_w[2] , \shft15_w[1] , \shft15_w[0] }), .shft14_w({
        \shft14_w[7] , \shft14_w[6] , \shft14_w[5] , \shft14_w[4] , 
        \shft14_w[3] , \shft14_w[2] , \shft14_w[1] , \shft14_w[0] }), 
        .fb_w_3(\fb_w[3] ), .fb_w_6(\fb_w[6] ), .fb_w_0(\fb_w[0] ), 
        .fb_w_7(\fb_w[7] ), .fb_w_1(\fb_w[1] ), .fb_w_2(\fb_w[2] ), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_566(N_566), .N_565(
        N_565), .N_568(N_568), .N_573(N_573));
    CFG3 #( .INIT(8'hCA) )  \codeOut_3[2]  (.A(\parity_w[2] ), .B(
        \dInp_reg_w[2] ), .C(datNotParity_w), .Y(\codeOut_3[2]_net_1 ));
    SLE \codeOut[5]  (.D(\codeOut_3[5]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(encoded[5]));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_165s_8s_0 tap_23 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft23_w({
        \shft23_w[7] , \shft23_w[6] , \shft23_w[5] , \shft23_w[4] , 
        \shft23_w[3] , \shft23_w[2] , \shft23_w[1] , \shft23_w[0] }), 
        .shft22_w({\shft22_w[7] , \shft22_w[6] , \shft22_w[5] , 
        \shft22_w[4] , \shft22_w[3] , \shft22_w[2] , \shft22_w[1] , 
        \shft22_w[0] }), .fb_w({\fb_w[7] , \fb_w[6] , \fb_w[5] , 
        \fb_w[4] , \fb_w[3] , \fb_w[2] , \fb_w[1] , \fb_w[0] }), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_574(N_574), .N_566(
        N_566), .N_568(N_568), .N_564(N_564), .N_570(N_570), .N_567(
        N_567), .N_565(N_565), .N_588(N_588));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_13s_8s_0 tap_26 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft26_w({
        \shft26_w[7] , \shft26_w[6] , \shft26_w[5] , \shft26_w[4] , 
        \shft26_w[3] , \shft26_w[2] , \shft26_w[1] , \shft26_w[0] }), 
        .fb_w({\fb_w[7] , \fb_w[6] , \fb_w[5] , \fb_w[4] , \fb_w[3] , 
        \fb_w[2] , \fb_w[1] , \fb_w[0] }), .shft25_w({\shft25_w[7] , 
        \shft25_w[6] , \shft25_w[5] , \shft25_w[4] , \shft25_w[3] , 
        \shft25_w[2] , \shft25_w[1] , \shft25_w[0] }), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_576(N_576), .N_583(
        N_583), .N_574(N_574), .N_572(N_572), .N_566(N_566), .N_575(
        N_575), .N_569(N_569));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_86s_8s_0 tap_13 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft13_w({
        \shft13_w[7] , \shft13_w[6] , \shft13_w[5] , \shft13_w[4] , 
        \shft13_w[3] , \shft13_w[2] , \shft13_w[1] , \shft13_w[0] }), 
        .shft12_w({\shft12_w[7] , \shft12_w[6] , \shft12_w[5] , 
        \shft12_w[4] , \shft12_w[3] , \shft12_w[2] , \shft12_w[1] , 
        \shft12_w[0] }), .fb_w({\fb_w[7] , \fb_w[6] , \fb_w[5] , 
        \fb_w[4] , \fb_w[3] , \fb_w[2] , \fb_w[1] }), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_568(N_568), .N_567(
        N_567), .N_574(N_574), .N_569(N_569), .N_576(N_576), .N_564(
        N_564), .N_565(N_565), .N_570(N_570), .N_575(N_575));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_113s_8s tap_16 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft16_w({\shft16_w[7] , 
        \shft16_w[6] , \shft16_w[5] , \shft16_w[4] , \shft16_w[3] , 
        \shft16_w[2] , \shft16_w[1] , \shft16_w[0] }), .shft15_w({
        \shft15_w[7] , \shft15_w[6] , \shft15_w[5] , \shft15_w[4] , 
        \shft15_w[3] , \shft15_w[2] , \shft15_w[1] , \shft15_w[0] }), 
        .fb_w_0(\fb_w[0] ), .fb_w_7(\fb_w[7] ), .fb_w_1(\fb_w[1] ), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_566(N_566), .N_567(
        N_567), .N_565(N_565), .N_574(N_574), .N_576(N_576), .N_583(
        N_583), .N_569(N_569), .N_564(N_564), .N_572(N_572), .N_568(
        N_568));
    CFG3 #( .INIT(8'hCA) )  \codeOut_3[5]  (.A(\parity_w[5] ), .B(
        \dInp_reg_w[5] ), .C(datNotParity_w), .Y(\codeOut_3[5]_net_1 ));
    CFG3 #( .INIT(8'hCA) )  \codeOut_3[4]  (.A(\parity_w[4] ), .B(
        \dInp_reg_w[4] ), .C(datNotParity_w), .Y(\codeOut_3[4]_net_1 ));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_42s_8s_0 tap_21 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft21_w({
        \shft21_w[7] , \shft21_w[6] , \shft21_w[5] , \shft21_w[4] , 
        \shft21_w[3] , \shft21_w[2] , \shft21_w[1] , \shft21_w[0] }), 
        .shft20_w({\shft20_w[7] , \shft20_w[6] , \shft20_w[5] , 
        \shft20_w[4] , \shft20_w[3] , \shft20_w[2] , \shft20_w[1] , 
        \shft20_w[0] }), .fb_w_1(\fb_w[3] ), .fb_w_3(\fb_w[5] ), 
        .fb_w_5(\fb_w[7] ), .fb_w_0(\fb_w[2] ), .fb_w_4(\fb_w[6] ), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_576(N_576), .N_564(
        N_564), .N_567(N_567), .N_565(N_565), .N_588(N_588), .N_570(
        N_570), .N_568(N_568), .N_575(N_575));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_42s_8s tap_11 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft11_w({\shft11_w[7] , 
        \shft11_w[6] , \shft11_w[5] , \shft11_w[4] , \shft11_w[3] , 
        \shft11_w[2] , \shft11_w[1] , \shft11_w[0] }), .shft10_w({
        \shft10_w[7] , \shft10_w[6] , \shft10_w[5] , \shft10_w[4] , 
        \shft10_w[3] , \shft10_w[2] , \shft10_w[1] , \shft10_w[0] }), 
        .fb_w_1(\fb_w[3] ), .fb_w_3(\fb_w[5] ), .fb_w_5(\fb_w[7] ), 
        .fb_w_0(\fb_w[2] ), .fb_w_4(\fb_w[6] ), .RSControl_0_NGRST(
        RSControl_0_NGRST), .N_576(N_576), .N_564(N_564), .N_567(N_567)
        , .N_565(N_565), .N_588(N_588), .N_570(N_570), .N_568(N_568), 
        .N_575(N_575));
    CFG2 #( .INIT(4'h6) )  \fb_w_i_o2[1]  (.A(\dInp_reg_w[1] ), .B(
        \pre_fb_w[1] ), .Y(\fb_w[1] ));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_127s_8s_0 tap_30 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft30_w({
        \shft30_w[7] , \shft30_w[6] , \shft30_w[5] , \shft30_w[4] , 
        \shft30_w[3] , \shft30_w[2] , \shft30_w[1] , \shft30_w[0] }), 
        .shft29_w({\shft29_w[7] , \shft29_w[6] , \shft29_w[5] , 
        \shft29_w[4] , \shft29_w[3] , \shft29_w[2] , \shft29_w[1] , 
        \shft29_w[0] }), .dInp_reg_w_3(\dInp_reg_w[6] ), .dInp_reg_w_2(
        \dInp_reg_w[5] ), .dInp_reg_w_0(\dInp_reg_w[3] ), .pre_fb_w_3(
        \pre_fb_w[6] ), .pre_fb_w_2(\pre_fb_w[5] ), .pre_fb_w_0(
        \pre_fb_w[3] ), .fb_w_4(\fb_w[4] ), .fb_w_7(\fb_w[7] ), 
        .fb_w_1(\fb_w[1] ), .fb_w_5(\fb_w[5] ), .fb_w_0(\fb_w[0] ), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_564(N_564), .N_570(
        N_570), .N_565(N_565), .N_567(N_567), .N_566(N_566), .N_569(
        N_569));
    SLE \codeOut[6]  (.D(\codeOut_3[6]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(encoded[6]));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_97s_8s_0 tap_24 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft24_w({
        \shft24_w[7] , \shft24_w[6] , \shft24_w[5] , \shft24_w[4] , 
        \shft24_w[3] , \shft24_w[2] , \shft24_w[1] , \shft24_w[0] }), 
        .shft23_w({\shft23_w[7] , \shft23_w[6] , \shft23_w[5] , 
        \shft23_w[4] , \shft23_w[3] , \shft23_w[2] , \shft23_w[1] , 
        \shft23_w[0] }), .fb_w({\fb_w[7] , \fb_w[6] , \fb_w[5] , 
        \fb_w[4] , \fb_w[3] , \fb_w[2] , \fb_w[1] , \fb_w[0] }), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_564(N_564), .N_567(
        N_567));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_171s_8s tap_14 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft14_w({\shft14_w[7] , 
        \shft14_w[6] , \shft14_w[5] , \shft14_w[4] , \shft14_w[3] , 
        \shft14_w[2] , \shft14_w[1] , \shft14_w[0] }), .shft13_w({
        \shft13_w[7] , \shft13_w[6] , \shft13_w[5] , \shft13_w[4] , 
        \shft13_w[3] , \shft13_w[2] , \shft13_w[1] , \shft13_w[0] }), 
        .fb_w_1(\fb_w[1] ), .fb_w_7(\fb_w[7] ), .fb_w_3(\fb_w[3] ), 
        .fb_w_5(\fb_w[5] ), .fb_w_0(\fb_w[0] ), .fb_w_6(\fb_w[6] ), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_583(N_583), .N_566(
        N_566), .N_569(N_569), .N_568(N_568), .N_572(N_572), .N_565(
        N_565), .N_567(N_567), .N_574(N_574));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_8s_8s_0 tap_22 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft22_w({\shft22_w[7] , 
        \shft22_w[6] , \shft22_w[5] , \shft22_w[4] , \shft22_w[3] , 
        \shft22_w[2] , \shft22_w[1] , \shft22_w[0] }), .shft21_w({
        \shft21_w[7] , \shft21_w[6] , \shft21_w[5] , \shft21_w[4] , 
        \shft21_w[3] , \shft21_w[2] , \shft21_w[1] , \shft21_w[0] }), 
        .fb_w_2(\fb_w[2] ), .fb_w_5(\fb_w[5] ), .fb_w_3(\fb_w[3] ), 
        .fb_w_6(\fb_w[6] ), .fb_w_0(\fb_w[0] ), .fb_w_7(\fb_w[7] ), 
        .fb_w_1(\fb_w[1] ), .RSControl_0_NGRST(RSControl_0_NGRST), 
        .N_566(N_566), .N_565(N_565));
    GND GND (.Y(GND_net_1));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_54s_8s tap_12 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft12_w({\shft12_w[7] , 
        \shft12_w[6] , \shft12_w[5] , \shft12_w[4] , \shft12_w[3] , 
        \shft12_w[2] , \shft12_w[1] , \shft12_w[0] }), .shft11_w({
        \shft11_w[7] , \shft11_w[6] , \shft11_w[5] , \shft11_w[4] , 
        \shft11_w[3] , \shft11_w[2] , \shft11_w[1] , \shft11_w[0] }), 
        .fb_w_5(\fb_w[5] ), .fb_w_2(\fb_w[2] ), .fb_w_0(\fb_w[0] ), 
        .fb_w_1(\fb_w[1] ), .fb_w_7(\fb_w[7] ), .RSControl_0_NGRST(
        RSControl_0_NGRST), .N_568(N_568), .N_575(N_575), .N_566(N_566)
        , .N_573(N_573), .N_567(N_567), .N_569(N_569), .N_572(N_572), 
        .N_565(N_565), .N_588(N_588));
    SLE \codeOut[3]  (.D(\codeOut_3[3]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(encoded[3]));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_30s_8s tap_5 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft5_w({\shft5_w[7] , \shft5_w[6] , 
        \shft5_w[5] , \shft5_w[4] , \shft5_w[3] , \shft5_w[2] , 
        \shft5_w[1] , \shft5_w[0] }), .shftOut_17_1({\shftOut_17_1[2] })
        , .shft4_w({\shft4_w[7] , \shft4_w[6] , \shft4_w[5] , 
        \shft4_w[4] , \shft4_w[3] , \shft4_w[2] , \shft4_w[1] , 
        \shft4_w[0] }), .fb_w_0(\fb_w[0] ), .fb_w_5(\fb_w[5] ), 
        .fb_w_3(\fb_w[3] ), .fb_w_6(\fb_w[6] ), .RSControl_0_NGRST(
        RSControl_0_NGRST), .N_566(N_566), .N_565(N_565), .N_572(N_572)
        , .N_575(N_575), .N_574(N_574), .N_564(N_564));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_127s_8s tap_2 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft2_w({\shft2_w[7] , \shft2_w[6] , 
        \shft2_w[5] , \shft2_w[4] , \shft2_w[3] , \shft2_w[2] , 
        \shft2_w[1] , \shft2_w[0] }), .shft1_w({\shft1_w[7] , 
        \shft1_w[6] , \shft1_w[5] , \shft1_w[4] , \shft1_w[3] , 
        \shft1_w[2] , \shft1_w[1] , \shft1_w[0] }), .fb_w_5(\fb_w[5] ), 
        .fb_w_0(\fb_w[0] ), .fb_w_1(\fb_w[1] ), .fb_w_4(\fb_w[4] ), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_567(N_567), .N_570(
        N_570), .N_565(N_565), .N_569(N_569), .N_566(N_566));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_91s_8s tap_1 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft1_w({\shft1_w[7] , \shft1_w[6] , 
        \shft1_w[5] , \shft1_w[4] , \shft1_w[3] , \shft1_w[2] , 
        \shft1_w[1] , \shft1_w[0] }), .shft0_w({\shft0_w[7] , 
        \shft0_w[6] , \shft0_w[5] , \shft0_w[4] , \shft0_w[3] , 
        \shft0_w[2] , \shft0_w[1] , \shft0_w[0] }), .fb_w_1(\fb_w[1] ), 
        .fb_w_5(\fb_w[5] ), .fb_w_3(\fb_w[3] ), .fb_w_0(\fb_w[0] ), 
        .fb_w_4(\fb_w[4] ), .RSControl_0_NGRST(RSControl_0_NGRST), 
        .N_564(N_564), .N_568(N_568), .N_572(N_572), .N_567(N_567), 
        .N_569(N_569));
    CFG2 #( .INIT(4'h6) )  \fb_w_i_o2[6]  (.A(\dInp_reg_w[6] ), .B(
        \pre_fb_w[6] ), .Y(\fb_w[6] ));
    CFG3 #( .INIT(8'hCA) )  \codeOut_3[1]  (.A(\parity_w[1] ), .B(
        \dInp_reg_w[1] ), .C(datNotParity_w), .Y(\codeOut_3[1]_net_1 ));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_16s_8s tap_4 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft4_w({\shft4_w[7] , \shft4_w[6] , 
        \shft4_w[5] , \shft4_w[4] , \shft4_w[3] , \shft4_w[2] , 
        \shft4_w[1] , \shft4_w[0] }), .shft3_w({\shft3_w[7] , 
        \shft3_w[6] , \shft3_w[5] , \shft3_w[4] , \shft3_w[3] , 
        \shft3_w[2] , \shft3_w[1] , \shft3_w[0] }), .fb_w_3(\fb_w[3] ), 
        .fb_w_4(\fb_w[4] ), .fb_w_2(\fb_w[2] ), .fb_w_6(\fb_w[6] ), 
        .fb_w_0(\fb_w[0] ), .fb_w_7(\fb_w[7] ), .fb_w_1(\fb_w[1] ), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_566(N_566), .N_565(
        N_565));
    CFG2 #( .INIT(4'h6) )  \fb_w_i_o2[2]  (.A(\dInp_reg_w[2] ), .B(
        \pre_fb_w[2] ), .Y(\fb_w[2] ));
    CFG2 #( .INIT(4'h6) )  \fb_w_i_o2[4]  (.A(\dInp_reg_w[4] ), .B(
        \pre_fb_w[4] ), .Y(\fb_w[4] ));
    CFG2 #( .INIT(4'h6) )  \fb_w_i_o2[5]  (.A(\dInp_reg_w[5] ), .B(
        \pre_fb_w[5] ), .Y(\fb_w[5] ));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_235s_8s tap_7 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft7_w({\shft7_w[7] , \shft7_w[6] , 
        \shft7_w[5] , \shft7_w[4] , \shft7_w[3] , \shft7_w[2] , 
        \shft7_w[1] , \shft7_w[0] }), .shft6_w({\shft6_w[7] , 
        \shft6_w[6] , \shft6_w[5] , \shft6_w[4] , \shft6_w[3] , 
        \shft6_w[2] , \shft6_w[1] , \shft6_w[0] }), .fb_w_1(\fb_w[1] ), 
        .fb_w_6(\fb_w[6] ), .fb_w_7(\fb_w[7] ), .fb_w_0(\fb_w[0] ), 
        .fb_w_3(\fb_w[3] ), .fb_w_5(\fb_w[5] ), .fb_w_4(\fb_w[4] ), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_564(N_564), .N_567(
        N_567));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_1s_8s tap_0 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft0_w({\shft0_w[7] , \shft0_w[6] , 
        \shft0_w[5] , \shft0_w[4] , \shft0_w[3] , \shft0_w[2] , 
        \shft0_w[1] , \shft0_w[0] }), .fb_w({\fb_w[7] , \fb_w[6] , 
        \fb_w[5] , \fb_w[4] , \fb_w[3] , \fb_w[2] , \fb_w[1] , 
        \fb_w[0] }), .RSControl_0_NGRST(RSControl_0_NGRST));
    CFG2 #( .INIT(4'h6) )  \fb_w_i_o2[7]  (.A(\dInp_reg_w[7] ), .B(
        \pre_fb_w[7] ), .Y(\fb_w[7] ));
    SLE \codeOut[1]  (.D(\codeOut_3[1]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(encoded[1]));
    CFG3 #( .INIT(8'hCA) )  \codeOut_3[0]  (.A(\parity_w[0] ), .B(
        \dInp_reg_w[0] ), .C(datNotParity_w), .Y(\codeOut_3[0]_net_1 ));
    CFG2 #( .INIT(4'h6) )  \fb_w_i_o2[0]  (.A(\dInp_reg_w[0] ), .B(
        \pre_fb_w[0] ), .Y(\fb_w[0] ));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_54s_8s_0 tap_20 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .shft20_w({
        \shft20_w[7] , \shft20_w[6] , \shft20_w[5] , \shft20_w[4] , 
        \shft20_w[3] , \shft20_w[2] , \shft20_w[1] , \shft20_w[0] }), 
        .shft19_w({\shft19_w[7] , \shft19_w[6] , \shft19_w[5] , 
        \shft19_w[4] , \shft19_w[3] , \shft19_w[2] , \shft19_w[1] , 
        \shft19_w[0] }), .fb_w_3(\fb_w[3] ), .fb_w_0(\fb_w[0] ), 
        .fb_w_5(\fb_w[5] ), .fb_w_2(\fb_w[2] ), .fb_w_1(\fb_w[1] ), 
        .fb_w_7(\fb_w[7] ), .RSControl_0_NGRST(RSControl_0_NGRST), 
        .N_588(N_588), .N_568(N_568), .N_575(N_575), .N_566(N_566), 
        .N_573(N_573), .N_567(N_567), .N_569(N_569), .N_572(N_572), 
        .N_565(N_565));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_8s_8s tap_10 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft10_w({\shft10_w[7] , 
        \shft10_w[6] , \shft10_w[5] , \shft10_w[4] , \shft10_w[3] , 
        \shft10_w[2] , \shft10_w[1] , \shft10_w[0] }), .shft9_w({
        \shft9_w[7] , \shft9_w[6] , \shft9_w[5] , \shft9_w[4] , 
        \shft9_w[3] , \shft9_w[2] , \shft9_w[1] , \shft9_w[0] }), 
        .fb_w_2(\fb_w[2] ), .fb_w_5(\fb_w[5] ), .fb_w_3(\fb_w[3] ), 
        .fb_w_6(\fb_w[6] ), .fb_w_0(\fb_w[0] ), .fb_w_7(\fb_w[7] ), 
        .fb_w_1(\fb_w[1] ), .RSControl_0_NGRST(RSControl_0_NGRST), 
        .N_566(N_566), .N_565(N_565));
    SLE \codeOut[0]  (.D(\codeOut_3[0]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(VCC_net_1), .ALn(
        RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(encoded[0]));
    TM_RSENC_TM_RSENC_0_rsEnc_lastTap_91s_8s tap_31 (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .dInp_reg_w({
        \dInp_reg_w[7] , \dInp_reg_w[6] , \dInp_reg_w[5] , 
        \dInp_reg_w[4] , \dInp_reg_w[3] , \dInp_reg_w[2] , 
        \dInp_reg_w[1] , \dInp_reg_w[0] }), .parity_w({\parity_w[7] , 
        \parity_w[6] , \parity_w[5] , \parity_w[4] , \parity_w[3] , 
        \parity_w[2] , \parity_w[1] , \parity_w[0] }), .pre_fb_w({
        \pre_fb_w[7] , \pre_fb_w[6] , \pre_fb_w[5] , \pre_fb_w[4] , 
        \pre_fb_w[3] , \pre_fb_w[2] , \pre_fb_w[1] , \pre_fb_w[0] }), 
        .conv_basis({conv_basis[7], conv_basis[6], conv_basis[5], 
        conv_basis[4], conv_basis[3], conv_basis[2], conv_basis[1], 
        conv_basis[0]}), .fb_w({\fb_w[7] , \fb_w[6] , \fb_w[5] , 
        \fb_w[4] , \fb_w[3] , \fb_w[2] , \fb_w[1] , \fb_w[0] }), 
        .shft30_w({\shft30_w[7] , \shft30_w[6] , \shft30_w[5] , 
        \shft30_w[4] , \shft30_w[3] , \shft30_w[2] , \shft30_w[1] , 
        \shft30_w[0] }), .RSControl_0_NGRST(RSControl_0_NGRST), 
        .hold0fb_w(hold0fb_w), .N_564(N_564), .N_569(N_569), .N_572(
        N_572), .N_568(N_568), .N_567(N_567));
    TM_RSENC_TM_RSENC_0_rsEnc_tap_13s_8s tap_6 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .shft6_w({\shft6_w[7] , \shft6_w[6] , 
        \shft6_w[5] , \shft6_w[4] , \shft6_w[3] , \shft6_w[2] , 
        \shft6_w[1] , \shft6_w[0] }), .shft5_w({\shft5_w[7] , 
        \shft5_w[6] , \shft5_w[5] , \shft5_w[4] , \shft5_w[3] , 
        \shft5_w[2] , \shft5_w[1] , \shft5_w[0] }), .fb_w_5(\fb_w[5] ), 
        .fb_w_3(\fb_w[3] ), .fb_w_2(\fb_w[2] ), .fb_w_7(\fb_w[7] ), 
        .fb_w_1(\fb_w[1] ), .fb_w_0(\fb_w[0] ), .fb_w_6(\fb_w[6] ), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .N_576(N_576), .N_583(
        N_583), .N_574(N_574), .N_566(N_566), .N_572(N_572), .N_575(
        N_575), .N_569(N_569));
    
endmodule


module TM_RSENC_TM_RSENC_0_tal1tab(
       Bit_Count_16dec_i_1,
       conv_basis,
       RSControl_0_DATAINP,
       RSControl_0_NGRST
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] conv_basis;
input  [7:0] RSControl_0_DATAINP;
input  RSControl_0_NGRST;

    wire VCC_net_1, \conv[4] , GND_net_1, \conv[5] , \conv[6] , 
        \conv[7] , \conv[0] , \conv[1] , \conv[2] , \conv[3] , N_24, 
        N_25;
    
    SLE \u[7]  (.D(\conv[7] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(conv_basis[7]));
    CFG2 #( .INIT(4'h6) )  \conv_i[1]  (.A(RSControl_0_DATAINP[5]), .B(
        RSControl_0_DATAINP[6]), .Y(\conv[1] ));
    CFG2 #( .INIT(4'h6) )  \conv_0_a2_0[2]  (.A(RSControl_0_DATAINP[0])
        , .B(RSControl_0_DATAINP[7]), .Y(N_24));
    SLE \u[5]  (.D(\conv[5] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(conv_basis[5]));
    CFG4 #( .INIT(16'h6996) )  \conv_0_a2[5]  (.A(
        RSControl_0_DATAINP[2]), .B(RSControl_0_DATAINP[3]), .C(N_25), 
        .D(RSControl_0_DATAINP[4]), .Y(\conv[5] ));
    SLE \u[4]  (.D(\conv[4] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(conv_basis[4]));
    SLE \u[0]  (.D(\conv[0] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(conv_basis[0]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \conv_0_a2[6]  (.A(
        RSControl_0_DATAINP[0]), .B(RSControl_0_DATAINP[6]), .C(
        \conv[4] ), .D(RSControl_0_DATAINP[7]), .Y(\conv[6] ));
    SLE \u[3]  (.D(\conv[3] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(conv_basis[3]));
    CFG3 #( .INIT(8'h96) )  \conv_0_a2[0]  (.A(RSControl_0_DATAINP[4]), 
        .B(RSControl_0_DATAINP[7]), .C(RSControl_0_DATAINP[2]), .Y(
        \conv[0] ));
    SLE \u[2]  (.D(\conv[2] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(conv_basis[2]));
    CFG3 #( .INIT(8'h96) )  \conv_0_a2[4]  (.A(RSControl_0_DATAINP[2]), 
        .B(RSControl_0_DATAINP[4]), .C(RSControl_0_DATAINP[3]), .Y(
        \conv[4] ));
    SLE \u[6]  (.D(\conv[6] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(conv_basis[6]));
    CFG2 #( .INIT(4'h6) )  \conv_0_a2_1[2]  (.A(RSControl_0_DATAINP[1])
        , .B(RSControl_0_DATAINP[5]), .Y(N_25));
    VCC VCC (.Y(VCC_net_1));
    SLE \u[1]  (.D(\conv[1] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(conv_basis[1]));
    CFG4 #( .INIT(16'h6996) )  \conv_0_a2[3]  (.A(
        RSControl_0_DATAINP[4]), .B(N_25), .C(RSControl_0_DATAINP[0]), 
        .D(RSControl_0_DATAINP[2]), .Y(\conv[3] ));
    CFG4 #( .INIT(16'h6996) )  \conv_0_a2[7]  (.A(
        RSControl_0_DATAINP[4]), .B(N_24), .C(RSControl_0_DATAINP[3]), 
        .D(RSControl_0_DATAINP[1]), .Y(\conv[7] ));
    CFG4 #( .INIT(16'h6996) )  \conv_0_a2[2]  (.A(
        RSControl_0_DATAINP[5]), .B(RSControl_0_DATAINP[1]), .C(N_24), 
        .D(RSControl_0_DATAINP[4]), .Y(\conv[2] ));
    
endmodule


module TM_RSENC_TM_RSENC_0_taltab(
       Bit_Count_16dec_i_1,
       TM_RSENC_0_CODEOUTP,
       encoded,
       RSControl_0_NGRST
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] TM_RSENC_0_CODEOUTP;
input  [7:0] encoded;
input  RSControl_0_NGRST;

    wire VCC_net_1, \dual[4] , GND_net_1, \dual[5] , \dual[6] , 
        \dual[7] , \dual[0] , \dual[1] , \dual[2] , \dual[3] , N_23, 
        \dual_0_a2_1[7]_net_1 ;
    
    SLE \z[4]  (.D(\dual[4] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TM_RSENC_0_CODEOUTP[4]));
    CFG4 #( .INIT(16'h6996) )  \dual_0_a2_1[7]  (.A(encoded[4]), .B(
        encoded[7]), .C(encoded[2]), .D(encoded[3]), .Y(
        \dual_0_a2_1[7]_net_1 ));
    SLE \z[3]  (.D(\dual[3] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TM_RSENC_0_CODEOUTP[3]));
    CFG4 #( .INIT(16'h6996) )  \dual_0_a2[1]  (.A(encoded[4]), .B(
        encoded[3]), .C(encoded[0]), .D(N_23), .Y(\dual[1] ));
    SLE \z[1]  (.D(\dual[1] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TM_RSENC_0_CODEOUTP[1]));
    GND GND (.Y(GND_net_1));
    SLE \z[2]  (.D(\dual[2] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TM_RSENC_0_CODEOUTP[2]));
    CFG4 #( .INIT(16'h6996) )  \dual_0_a2[6]  (.A(encoded[6]), .B(
        encoded[5]), .C(encoded[3]), .D(encoded[0]), .Y(\dual[6] ));
    CFG4 #( .INIT(16'h6996) )  \dual_0_a2[0]  (.A(encoded[7]), .B(
        encoded[2]), .C(encoded[0]), .D(N_23), .Y(\dual[0] ));
    CFG3 #( .INIT(8'h96) )  \dual_0_a2[3]  (.A(encoded[7]), .B(
        encoded[2]), .C(\dual[5] ), .Y(\dual[3] ));
    CFG4 #( .INIT(16'h6996) )  \dual_0_a2[2]  (.A(encoded[7]), .B(
        encoded[4]), .C(N_23), .D(encoded[5]), .Y(\dual[2] ));
    CFG3 #( .INIT(8'h96) )  \dual_0_a2[7]  (.A(\dual_0_a2_1[7]_net_1 ), 
        .B(encoded[5]), .C(N_23), .Y(\dual[7] ));
    CFG4 #( .INIT(16'h6996) )  \dual_0_a2[5]  (.A(encoded[5]), .B(
        encoded[3]), .C(encoded[0]), .D(N_23), .Y(\dual[5] ));
    VCC VCC (.Y(VCC_net_1));
    SLE \z[6]  (.D(\dual[6] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TM_RSENC_0_CODEOUTP[6]));
    SLE \z[5]  (.D(\dual[5] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TM_RSENC_0_CODEOUTP[5]));
    CFG2 #( .INIT(4'h6) )  \dual_0_a2_0[0]  (.A(encoded[6]), .B(
        encoded[1]), .Y(N_23));
    SLE \z[0]  (.D(\dual[0] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TM_RSENC_0_CODEOUTP[0]));
    CFG3 #( .INIT(8'h96) )  \dual_0_a2[4]  (.A(encoded[3]), .B(
        encoded[0]), .C(encoded[2]), .Y(\dual[4] ));
    SLE \z[7]  (.D(\dual[7] ), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(RSControl_0_NGRST), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TM_RSENC_0_CODEOUTP[7]));
    
endmodule


module TM_RSENC_TM_RSENC_0_CORERSENC_16s_255s_8s_1s_1s_19s_223s(
       Bit_Count_16dec_i_1,
       RSControl_0_DATAINP,
       TM_RSENC_0_CODEOUTP,
       TM_RSENC_0_RFD,
       RSControl_0_NGRST,
       TM_RSENC_0_RFS,
       RSControl_0_START,
       TM_RSENC_0_RDY
    );
input  [3:3] Bit_Count_16dec_i_1;
input  [7:0] RSControl_0_DATAINP;
output [7:0] TM_RSENC_0_CODEOUTP;
output TM_RSENC_0_RFD;
input  RSControl_0_NGRST;
output TM_RSENC_0_RFS;
input  RSControl_0_START;
output TM_RSENC_0_RDY;

    wire hold0fb_w, datNotParity_w, \conv_basis[0] , \conv_basis[1] , 
        \conv_basis[2] , \conv_basis[3] , \conv_basis[4] , 
        \conv_basis[5] , \conv_basis[6] , \conv_basis[7] , 
        \encoded[0] , \encoded[1] , \encoded[2] , \encoded[3] , 
        \encoded[4] , \encoded[5] , \encoded[6] , \encoded[7] , 
        GND_net_1, VCC_net_1;
    
    TM_RSENC_TM_RSENC_0_rsEnc_SM_223s_16s_255s_8s_1s_1s_4s 
        TM_RSENC_TM_RSENC_0_rsEnc_SM_0 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .hold0fb_w(hold0fb_w), 
        .TM_RSENC_0_RFD(TM_RSENC_0_RFD), .RSControl_0_NGRST(
        RSControl_0_NGRST), .TM_RSENC_0_RFS(TM_RSENC_0_RFS), 
        .datNotParity_w(datNotParity_w), .RSControl_0_START(
        RSControl_0_START), .TM_RSENC_0_RDY(TM_RSENC_0_RDY));
    VCC VCC (.Y(VCC_net_1));
    TM_RSENC_TM_RSENC_0_gfIIR_8s gfIIR_0 (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .encoded({\encoded[7] , \encoded[6] , 
        \encoded[5] , \encoded[4] , \encoded[3] , \encoded[2] , 
        \encoded[1] , \encoded[0] }), .conv_basis({\conv_basis[7] , 
        \conv_basis[6] , \conv_basis[5] , \conv_basis[4] , 
        \conv_basis[3] , \conv_basis[2] , \conv_basis[1] , 
        \conv_basis[0] }), .RSControl_0_NGRST(RSControl_0_NGRST), 
        .datNotParity_w(datNotParity_w), .hold0fb_w(hold0fb_w));
    TM_RSENC_TM_RSENC_0_tal1tab \convert_inp.tal1tab_0  (
        .Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), .conv_basis({
        \conv_basis[7] , \conv_basis[6] , \conv_basis[5] , 
        \conv_basis[4] , \conv_basis[3] , \conv_basis[2] , 
        \conv_basis[1] , \conv_basis[0] }), .RSControl_0_DATAINP({
        RSControl_0_DATAINP[7], RSControl_0_DATAINP[6], 
        RSControl_0_DATAINP[5], RSControl_0_DATAINP[4], 
        RSControl_0_DATAINP[3], RSControl_0_DATAINP[2], 
        RSControl_0_DATAINP[1], RSControl_0_DATAINP[0]}), 
        .RSControl_0_NGRST(RSControl_0_NGRST));
    GND GND (.Y(GND_net_1));
    TM_RSENC_TM_RSENC_0_taltab \ccsds.taltab_0  (.Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .TM_RSENC_0_CODEOUTP({
        TM_RSENC_0_CODEOUTP[7], TM_RSENC_0_CODEOUTP[6], 
        TM_RSENC_0_CODEOUTP[5], TM_RSENC_0_CODEOUTP[4], 
        TM_RSENC_0_CODEOUTP[3], TM_RSENC_0_CODEOUTP[2], 
        TM_RSENC_0_CODEOUTP[1], TM_RSENC_0_CODEOUTP[0]}), .encoded({
        \encoded[7] , \encoded[6] , \encoded[5] , \encoded[4] , 
        \encoded[3] , \encoded[2] , \encoded[1] , \encoded[0] }), 
        .RSControl_0_NGRST(RSControl_0_NGRST));
    
endmodule


module TM_RSENC(
       Bit_Count_16dec_i_1,
       RSControl_0_DATAINP,
       TM_RSENC_0_CODEOUTP,
       TM_RSENC_0_RFD,
       RSControl_0_NGRST,
       TM_RSENC_0_RFS,
       RSControl_0_START,
       TM_RSENC_0_RDY
    );
input  [3:3] Bit_Count_16dec_i_1;
input  [7:0] RSControl_0_DATAINP;
output [7:0] TM_RSENC_0_CODEOUTP;
output TM_RSENC_0_RFD;
input  RSControl_0_NGRST;
output TM_RSENC_0_RFS;
input  RSControl_0_START;
output TM_RSENC_0_RDY;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    TM_RSENC_TM_RSENC_0_CORERSENC_16s_255s_8s_1s_1s_19s_223s 
        TM_RSENC_0 (.Bit_Count_16dec_i_1({Bit_Count_16dec_i_1[3]}), 
        .RSControl_0_DATAINP({RSControl_0_DATAINP[7], 
        RSControl_0_DATAINP[6], RSControl_0_DATAINP[5], 
        RSControl_0_DATAINP[4], RSControl_0_DATAINP[3], 
        RSControl_0_DATAINP[2], RSControl_0_DATAINP[1], 
        RSControl_0_DATAINP[0]}), .TM_RSENC_0_CODEOUTP({
        TM_RSENC_0_CODEOUTP[7], TM_RSENC_0_CODEOUTP[6], 
        TM_RSENC_0_CODEOUTP[5], TM_RSENC_0_CODEOUTP[4], 
        TM_RSENC_0_CODEOUTP[3], TM_RSENC_0_CODEOUTP[2], 
        TM_RSENC_0_CODEOUTP[1], TM_RSENC_0_CODEOUTP[0]}), 
        .TM_RSENC_0_RFD(TM_RSENC_0_RFD), .RSControl_0_NGRST(
        RSControl_0_NGRST), .TM_RSENC_0_RFS(TM_RSENC_0_RFS), 
        .RSControl_0_START(RSControl_0_START), .TM_RSENC_0_RDY(
        TM_RSENC_0_RDY));
    
endmodule


module Glue_Logic_Z10(
       Glue_Logic_0_USER_RA_TRP1_1,
       Glue_Logic_0_MSG_WA_TRP1,
       CoreAPB3_0_APBmslave3_PRDATA,
       Glue_Logic_0_MSG_TRP1,
       Glue_Logic_0_Flag_Int_0,
       CoreAPB3_0_APBmslave3_PADDR,
       CoreAPB3_0_APBmslave3_PWDATA,
       CPU_W_HDL_R_0_TM_Packet_Counter,
       CLTU_0_TC_Packet_Counter,
       CLTU_0_TC_Error_Counter,
       COREEDAC_1_DATA_OUT,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       OSC_0_XTLOSC_O2F,
       Glue_Logic_0_USER_REN_TRP1,
       Glue_Logic_0_Flag_B_Tx,
       Glue_Logic_0_Flag_B_Rx,
       TXD4_net_0,
       Flag_RX,
       Glue_Logic_0_USER_WEN_TRP1,
       CoreAPB3_0_APBmslave3_PREADY,
       HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish,
       CPU_W_HDL_R_0_Flag_A_Tx_Finish,
       HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish,
       CPU_W_HDL_R_0_Flag_B_Tx_Finish,
       CoreAPB3_0_APBmslave3_PWRITE,
       Switch_0_EnOut,
       CLTU_0_Flag_RX_ing,
       test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx,
       CoreAPB3_0_APBmslave3_PENABLE,
       iPSELS_raw23
    );
output [3:0] Glue_Logic_0_USER_RA_TRP1_1;
output [9:0] Glue_Logic_0_MSG_WA_TRP1;
output [31:0] CoreAPB3_0_APBmslave3_PRDATA;
output [7:0] Glue_Logic_0_MSG_TRP1;
output [0:0] Glue_Logic_0_Flag_Int_0;
input  [31:0] CoreAPB3_0_APBmslave3_PADDR;
input  [31:0] CoreAPB3_0_APBmslave3_PWDATA;
input  [31:0] CPU_W_HDL_R_0_TM_Packet_Counter;
input  [31:0] CLTU_0_TC_Packet_Counter;
input  [31:0] CLTU_0_TC_Error_Counter;
input  [31:0] COREEDAC_1_DATA_OUT;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  OSC_0_XTLOSC_O2F;
output Glue_Logic_0_USER_REN_TRP1;
output Glue_Logic_0_Flag_B_Tx;
output Glue_Logic_0_Flag_B_Rx;
output TXD4_net_0;
output Flag_RX;
output Glue_Logic_0_USER_WEN_TRP1;
output CoreAPB3_0_APBmslave3_PREADY;
input  HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish;
input  CPU_W_HDL_R_0_Flag_A_Tx_Finish;
input  HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish;
input  CPU_W_HDL_R_0_Flag_B_Tx_Finish;
input  CoreAPB3_0_APBmslave3_PWRITE;
input  Switch_0_EnOut;
input  CLTU_0_Flag_RX_ing;
input  test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx;
input  CoreAPB3_0_APBmslave3_PENABLE;
input  iPSELS_raw23;

    wire Flag_Enable_net_1, Flag_Enable_i_0, \APB_ADDRESS[27]_net_1 , 
        VCC_net_1, GND_net_1, \APB_ADDRESS[28]_net_1 , 
        \APB_ADDRESS[29]_net_1 , \APB_ADDRESS[30]_net_1 , 
        \APB_ADDRESS[31]_net_1 , \APB_ADDRESS[12]_net_1 , 
        \APB_ADDRESS[13]_net_1 , \APB_ADDRESS[14]_net_1 , 
        \APB_ADDRESS[15]_net_1 , \APB_ADDRESS[16]_net_1 , 
        \APB_ADDRESS[17]_net_1 , \APB_ADDRESS[18]_net_1 , 
        \APB_ADDRESS[19]_net_1 , \APB_ADDRESS[20]_net_1 , 
        \APB_ADDRESS[21]_net_1 , \APB_ADDRESS[22]_net_1 , 
        \APB_ADDRESS[23]_net_1 , \APB_ADDRESS[24]_net_1 , 
        \APB_ADDRESS[25]_net_1 , \APB_ADDRESS[26]_net_1 , 
        \APB_ADDRESS[2]_net_1 , Flag_Enable_1_sqmuxa, 
        \APB_ADDRESS[3]_net_1 , \APB_ADDRESS[4]_net_1 , N_49_i, 
        \Byte_Count[0]_net_1 , N_145_i_0, \Byte_Count[1]_net_1 , 
        N_1029_i_0, \APB_ADDRESS[5]_net_1 , \APB_ADDRESS[10]_net_1 , 
        \APB_ADDRESS[11]_net_1 , \PRDATA_14[27] , un1_PRDATA47_1_i_0, 
        \PRDATA_14[28] , \PRDATA_14[29] , \PRDATA_14[30] , 
        \PRDATA_14[31] , un1_PADDR_1_cry_0_Y, N_986_i_0, 
        un1_PADDR_1_cry_1_S, un1_PADDR_1_cry_2_S, un1_PADDR_1_cry_3_S, 
        un1_PADDR_1_cry_4_S, un1_PADDR_1_cry_5_S, un1_PADDR_1_cry_6_S, 
        un1_PADDR_1_cry_7_S, un1_PADDR_1_cry_8_S, un1_PADDR_1_s_9_S, 
        \PRDATA_14[12] , \PRDATA_14[13] , \PRDATA_14[14] , 
        \PRDATA_14[15] , \PRDATA_14[16] , \PRDATA_14[17] , 
        \PRDATA_14[18] , \PRDATA_14[19] , \PRDATA_14[20] , 
        \PRDATA_14[21] , \PRDATA_14[22] , \PRDATA_14[23] , 
        \PRDATA_14[24] , \PRDATA_14[25] , \PRDATA_14[26] , 
        \MSG_TRP1_13[5] , \MSG_TRP1_13[6] , N_990, \PRDATA_14[0] , 
        \PRDATA_14[1] , \PRDATA_14[2] , \PRDATA_14[3] , 
        PRDATA_N_5_mux_0_i_0, \PRDATA_14[5] , \PRDATA_14[6] , 
        \PRDATA_14[7] , \PRDATA_14[8] , \PRDATA_14[9] , 
        \PRDATA_14[10] , \PRDATA_14[11] , N_994, N_993, N_992, N_991, 
        \MSG_TRP1_13[4] , USER_REN_TRP1ce_net_1, 
        un1_Flag_Int_1_sqmuxa_1, Flag_Int_1_sqmuxa_1_i_0_0_net_1, 
        Flag_B_Tx18_net_1, Flag_B_Tx_0_sqmuxa_1_i_0, Flag_B_Rx18_net_1, 
        Flag_B_Rx_0_sqmuxa_1_i_0_0_net_1, Flag_A_Tx18_net_1, 
        Flag_A_Tx_0_sqmuxa_1_i_0, Flag_A_Rx18_net_1, 
        Flag_A_Rx_0_sqmuxa_1_i_0_0_net_1, Flag_Enable1_net_1, 
        Flag_Enable1_1_sqmuxa_1, Flag_Enable1_1_sqmuxa_2_i_0_net_1, 
        Flag_Enable_1_sqmuxa_1_i_0_net_1, PREADY_9, 
        pos1_Flag_A_HDL_Rec_Finish_net_1, pos1_Flag_A_Tx_Finish_net_1, 
        pos1_Flag_B_HDL_Rec_Finish_net_1, pos1_Flag_B_Tx_Finish_net_1, 
        pos2_Flag_A_HDL_Rec_Finish_net_1, pos2_Flag_A_Tx_Finish_net_1, 
        pos2_Flag_B_HDL_Rec_Finish_net_1, pos2_Flag_B_Tx_Finish_net_1, 
        un1_PADDR_1_cry_0_net_1, N_984, un1_PADDR_1_cry_1_net_1, 
        un1_PADDR_1_cry_2_net_1, un1_PADDR_1_cry_3_net_1, 
        un1_PADDR_1_cry_4_net_1, un1_PADDR_1_cry_5_net_1, 
        un1_PADDR_1_cry_6_net_1, un1_PADDR_1_cry_7_net_1, N_982, 
        un25_TXB_0_a2_0_net_1, N_980, un1_PADDR_1_cry_8_net_1, 
        Flag_Int_1_sqmuxa_1_i_0_0_1_0_net_1, PRDATA30_2_0_1_net_1, 
        PRDATA30_2_0_sx_6_net_1, PRDATA30_2_0_sx_4_net_1, 
        PRDATA30_2_0_sx_5_net_1, PRDATA34_2_0, PRDATA30_2_0_sx_net_1, 
        un1_PRDATA30_4_0_a3_0_4_sx_net_1, PRDATA30_2_0_x_0_net_1, 
        un1_PRDATA30_4_0_a3_0_4_x_net_1, un1_m2_e_2_2_1, PRDATA30_26_3, 
        un1_PRDATA30_4_0_a3_0_sx_0_net_1, un1_PRDATA30_4_0_a3_0_1, 
        PRDATA30_26_4, un1_PRDATA30_4_0_i_a2_1_0_net_1, 
        un1_PRDATA30_4_0_i_a2_sx_net_1, N_629, PRDATA30_2_0_sx_2_net_1, 
        PRDATA30_2_0_sx_3_net_1, PRDATA30_2_0_2_net_1, 
        PRDATA37_0_net_1, PRDATA37_2_sx_net_1, PRDATA37_2_net_1, 
        un1_PRDATA30_4_0_a3_0_3, PRDATA30_2_0_3_RNIUOJ6_net_1, N_1406, 
        un1_PRDATA47_1_i_0_a2_N_3L3_1, PRDATA38_1_0_net_1, 
        un1_PRDATA47_1_i_0_a2_1, \APB_ADDRESS_RNI3P7M[13]_net_1 , 
        N_506, g2_8_net_1, PRDATA36_1_net_1, PRDATA36_2_net_1, 
        PRDATA37_1_0, g0_sx, g0_1_net_1, un1_m2_e_2_2_1_0, 
        PRDATA38_1_0_0_net_1, N_1025, PRDATA30_2_0_3_net_1, 
        PRDATA30_2_0_4_net_1, \PRDATA_14_iv_0_2_sx[8]_net_1 , 
        \PRDATA_14_iv_0_2_0[8]_net_1 , N_510, 
        \PRDATA_14_iv_0_2[8]_net_1 , PRDATA36_3_net_1, 
        \PRDATA_14_iv_0_1[3]_net_1 , \PRDATA_14_iv_0[3]_net_1 , 
        PRDATA30_2_0_x_net_1, un1_PRDATA30_4_0_o3_sx_0, 
        un1_PRDATA30_4_0_o3_4_0, N_660, Flag_m3_e_1_1, 
        un1_PRDATA30_4_0_o3_sx, PRDATA_m2_0, 
        \PRDATA_14_0_iv_0_sx_sx[9]_net_1 , 
        \PRDATA_14_0_iv_0_sx[9]_net_1 , PRDATA30_2_0_sx_0_net_1, 
        un1_PRDATA30_4_0_o3_4_0_sx, un1_PRDATA30_4_0_a3_0, N_658, 
        N_651, \PRDATA_14_iv_2[5]_net_1 , \PRDATA_14_iv_sx[5]_net_1 , 
        un1_PRDATA39_1, un1_PRDATA30_4_0_o3_4, un1_m2_e_2, 
        \PRDATA_14_iv_2[6]_net_1 , \PRDATA_14_iv_sx[6]_net_1 , 
        \PRDATA_14_iv_0_sx[7]_net_1 , \PRDATA_14_iv_0_2[7]_net_1 , 
        \PRDATA_14_iv_2[3]_net_1 , \PRDATA_14_iv_sx[3]_net_1 , 
        \PRDATA_14_iv_0_o2_0_0[4]_net_1 , 
        \PRDATA_14_iv_0_o2_0_x_RNO[4]_net_1 , 
        \PRDATA_14_iv_0_o2_0_x[4]_net_1 , PRDATA33_0_net_1, 
        PRDATA33_3_x_net_1, Flag_m3_e_1_1_1, 
        un1_PRDATA30_4_0_o3_4_sx_sx_0_net_1, 
        un1_PRDATA30_4_0_o3_4_1_sx_sx_net_1, un1_PRDATA30_4_0_o3_4_1_0, 
        \PRDATA_14_iv_0_3_RNO[8]_net_1 , \PRDATA_14_iv_0_3[8]_net_1 , 
        PRDATA33_net_1, PRDATA33_1_0_0_o2_x_net_1, 
        PRDATA33_1_0_0_o2_1_net_1, PRDATA33_4_net_1, 
        \PRDATA_14_iv_0_o2_1_1[4]_net_1 , un1_PRDATA30_4_0_o3_4_2, 
        \PRDATA_14_iv_1_1[0]_net_1 , \PRDATA_14_iv_1_sx[0]_net_1 , 
        \PRDATA_14_iv_1[0]_net_1 , un1_m2_e_0_1_sx, un1_m2_e_0_1, 
        N_507, \PRDATA_14_0_iv_0_sx[10]_net_1 , 
        \PRDATA_14_0_iv_0_1[10]_net_1 , \PRDATA_14_0_iv_0_1[9]_net_1 , 
        un25_TXB_0_o2_0_x_net_1, PRDATA33_6_net_1, 
        un25_TXB_0_o2_0_3_net_1, un25_TXB_0_o2_0_0_net_1, 
        un25_TXB_0_o2_0_1_net_1, un25_TXB_0_o2_0_2_net_1, 
        un1_PRDATA30_4_0_o3_0, \PRDATA_14_iv_0_1_1_0[7]_net_1 , 
        \PRDATA_14_iv_0_1[7] , N_977, Flag_Enable_RNIDIIB1_net_1, 
        Flag_m3_e_1, g0_1_0_net_1, g0_3_3_net_1, PRDATA32_4, 
        g2_6_net_1, g2_5_net_1, g0_3_4_net_1, PRDATA34_26, 
        PRDATA30_2_0_RNIUQLC2_net_1, PRDATA30_1_0_0_a3_0_net_1, 
        PRDATA35_1_0_0_a3_RNIV4QV_net_1, N_502, 
        \PRDATA_14_iv_0_o2_1_RNI894C2[4]_net_1 , 
        un1_PRDATA47_1_i_0_a2_0, \PRDATA_14_iv_2_1[5]_net_1 , 
        \PRDATA_14_iv_0[5]_net_1 , PRDATA30, \PRDATA_14_iv_0[6]_net_1 , 
        \PRDATA_14_iv_2_1[6]_net_1 , PRDATA_m2_0_a2_2, 
        PRDATA_N_5_mux_0_i_1_net_1, PRDATA_m2_0_a2_0, 
        USER_REN_TRP1ce_1_net_1, \PRDATA_14_0_iv_1_1[20]_net_1 , 
        \PRDATA_14_0_iv_1[20]_net_1 , \PRDATA_14_0_iv_1_1[25]_net_1 , 
        \PRDATA_14_0_iv_1[25]_net_1 , \PRDATA_14_0_iv_1_1[12]_net_1 , 
        \PRDATA_14_0_iv_1[12]_net_1 , \PRDATA_14_0_iv_0_1_1[27]_net_1 , 
        \PRDATA_14_0_iv_0_1[27]_net_1 , \PRDATA_14_0_iv_1_1[11]_net_1 , 
        \PRDATA_14_0_iv_1[11]_net_1 , \PRDATA_14_0_iv_1_1[19]_net_1 , 
        \PRDATA_14_0_iv_1[19]_net_1 , \PRDATA_14_0_iv_0_1_1[28]_net_1 , 
        \PRDATA_14_0_iv_0_1[28]_net_1 , \PRDATA_14_0_iv_1_1[22]_net_1 , 
        \PRDATA_14_0_iv_1[22]_net_1 , \PRDATA_14_0_iv_0_1_1[26]_net_1 , 
        \PRDATA_14_0_iv_0_1[26]_net_1 , 
        \PRDATA_14_0_iv_0_1_1[24]_net_1 , 
        \PRDATA_14_0_iv_0_1[24]_net_1 , 
        \PRDATA_14_0_iv_0_1_1[21]_net_1 , 
        \PRDATA_14_0_iv_0_1[21]_net_1 , \PRDATA_14_0_iv_1_1[13]_net_1 , 
        \PRDATA_14_0_iv_1[13]_net_1 , \PRDATA_14_0_iv_0_1_1[29]_net_1 , 
        \PRDATA_14_0_iv_0_1[29]_net_1 , 
        \PRDATA_14_0_iv_0_1_1[16]_net_1 , 
        \PRDATA_14_0_iv_0_1[16]_net_1 , \MSG_TRP1_13_3_i_m2_1_1[3] , 
        \MSG_TRP1_13_3_1_1[6] , \MSG_TRP1_13_3_1_1[5] , 
        \MSG_TRP1_13_3_i_m2_1_1[7] , \MSG_TRP1_13_3_i_m2_1_1[2] , 
        \MSG_TRP1_13_3_i_m2_1_1[0] , \MSG_TRP1_13_3_i_m2_1_1[1] , 
        \MSG_TRP1_13_3_1_1[4] , Flag_Enable1_1_sqmuxa_1_1, 
        PRDATA_m1_0_a2_0, PRDATA33_3_net_1, PRDATA35_1_0_0_a3_1_net_1, 
        un1_PRDATA30_4_0_o3_0_13, un1_PRDATA30_4_0_o3_0_12, 
        un1_PRDATA30_4_0_o3_0_11, un1_PRDATA30_4_0_o3_0_10, N_644, 
        un1_PRDATA30_4_0_o3_0_14, N_138, N_1000, N_985, 
        PRDATA_m1_0_a2_2, \TM_Packet_Counter_m[31] , 
        \TM_Packet_Counter_m[15] , \TC_Packet_Counter_m[3] , N_618, 
        N_536, N_528, \TC_Error_Counter_m[6] , 
        \TM_Packet_Counter_m[17] , N_524, \TM_Packet_Counter_m[2] , 
        \TC_Error_Counter_m[2] , \TC_Error_Counter_m[5] , 
        \TM_Packet_Counter_m[1] , \TC_Error_Counter_m[1] , N_563, 
        \TM_Packet_Counter_m[23] , N_540, 
        \PRDATA_14_0_iv_0_0[10]_net_1 , \PRDATA_14_0_iv_0_0[9]_net_1 , 
        \PRDATA_14_iv_0[1]_net_1 , \PRDATA_14_iv_0[31]_net_1 , 
        \PRDATA_14_0_iv_0[17]_net_1 , \PRDATA_14_0_iv_0_0[18]_net_1 , 
        \PRDATA_14_0_iv_0_0[30]_net_1 , \PRDATA_14_0_iv_0_0[14]_net_1 , 
        \PRDATA_14_iv_0[2]_net_1 , \PRDATA_14_0_iv_0[15]_net_1 , 
        \PRDATA_14_0_iv_0[23]_net_1 , PREADY_9_0_0_tz_net_1, 
        Flag_Int_0_sqmuxa_2_net_1, \PRDATA_14_0_iv_1[17]_net_1 , 
        \PRDATA_14_0_iv_0_1[18]_net_1 , \PRDATA_14_0_iv_0_1[30]_net_1 , 
        \PRDATA_14_0_iv_0_1[14]_net_1 , \PRDATA_14_0_iv_1[15]_net_1 , 
        \PRDATA_14_0_iv_1[23]_net_1 , un1_m2_e_1, 
        \PRDATA_14_iv_2[0]_net_1 , \PRDATA_14_iv_2[1]_net_1 , 
        \PRDATA_14_iv_2[31]_net_1 , \PRDATA_14_iv_2[2]_net_1 , 
        un1_PRDATA47_1_i_0_a2_1_0, Flag_m1_e_1, un1_N_5_mux_2, 
        un1_N_5_mux_0_0;
    
    CFG2 #( .INIT(4'h1) )  PREADY_9_0_o2_RNIO2EL1 (.A(N_984), .B(N_985)
        , .Y(N_986_i_0));
    SLE \MSG_WA_TRP1[8]  (.D(un1_PADDR_1_cry_8_S), .CLK(
        OSC_0_XTLOSC_O2F), .EN(N_986_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_MSG_WA_TRP1[8]));
    SLE \USER_RA_TRP1[1]  (.D(\APB_ADDRESS[3]_net_1 ), .CLK(
        OSC_0_XTLOSC_O2F), .EN(Flag_Enable_1_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_USER_RA_TRP1_1[1]));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_iv_0[7]  (.A(
        COREEDAC_1_DATA_OUT[31]), .B(\PRDATA_14_iv_0_sx[7]_net_1 ), .C(
        \PRDATA_14_iv_0_2[7]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[7] ));
    CFG4 #( .INIT(16'h8000) )  PRDATA36_3 (.A(PRDATA36_1_net_1), .B(
        PRDATA30_26_3), .C(PRDATA36_2_net_1), .D(PRDATA30_26_4), .Y(
        PRDATA36_3_net_1));
    SLE pos1_Flag_B_Tx_Finish (.D(CPU_W_HDL_R_0_Flag_B_Tx_Finish), 
        .CLK(OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pos1_Flag_B_Tx_Finish_net_1));
    SLE Flag_Enable (.D(Flag_Enable_1_sqmuxa), .CLK(OSC_0_XTLOSC_O2F), 
        .EN(Flag_Enable_1_sqmuxa_1_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Flag_Enable_net_1));
    CFG4 #( .INIT(16'h2000) )  un1_PRDATA47_1_i_0_a2_0_0 (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        CoreAPB3_0_APBmslave3_PWRITE), .C(
        CoreAPB3_0_APBmslave3_PENABLE), .D(iPSELS_raw23), .Y(
        un1_PRDATA47_1_i_0_a2_0));
    SLE \PRDATA[5]  (.D(\PRDATA_14[5] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[5]));
    SLE \PRDATA[30]  (.D(\PRDATA_14[30] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[30]));
    ARI1 #( .INIT(20'h4AA00) )  un1_PADDR_1_cry_5 (.A(VCC_net_1), .B(
        CoreAPB3_0_APBmslave3_PADDR[5]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un1_PADDR_1_cry_4_net_1), .S(un1_PADDR_1_cry_5_S), .Y(), 
        .FCO(un1_PADDR_1_cry_5_net_1));
    CFG4 #( .INIT(16'hFFFE) )  PRDATA30_2_0_sx_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[21]), .B(
        CoreAPB3_0_APBmslave3_PADDR[26]), .C(
        CoreAPB3_0_APBmslave3_PADDR[20]), .D(
        CoreAPB3_0_APBmslave3_PADDR[27]), .Y(PRDATA30_2_0_sx_0_net_1));
    CFG4 #( .INIT(16'hEAC0) )  Flag_Int_1_sqmuxa_1_i_0_0_1_0 (.A(
        CPU_W_HDL_R_0_Flag_B_Tx_Finish), .B(
        CPU_W_HDL_R_0_Flag_A_Tx_Finish), .C(TXD4_net_0), .D(
        Glue_Logic_0_Flag_B_Tx), .Y(
        Flag_Int_1_sqmuxa_1_i_0_0_1_0_net_1));
    CFG4 #( .INIT(16'hFDDD) )  \PRDATA_14_iv_2[5]  (.A(
        \PRDATA_14_iv_2_1[5]_net_1 ), .B(\PRDATA_14_iv_0[5]_net_1 ), 
        .C(Switch_0_EnOut), .D(PRDATA30), .Y(\PRDATA_14_iv_2[5]_net_1 )
        );
    CFG4 #( .INIT(16'h80CC) )  \PRDATA_14_iv_0_1_0[7]  (.A(
        CLTU_0_TC_Error_Counter[7]), .B(PRDATA34_2_0), .C(
        PRDATA38_1_0_net_1), .D(\PRDATA_14_iv_0_1_1_0[7]_net_1 ), .Y(
        \PRDATA_14_iv_0_1[7] ));
    CFG4 #( .INIT(16'h4657) )  \MSG_TRP1_RNO_0[6]  (.A(
        \Byte_Count[1]_net_1 ), .B(\Byte_Count[0]_net_1 ), .C(
        CoreAPB3_0_APBmslave3_PWDATA[22]), .D(
        CoreAPB3_0_APBmslave3_PWDATA[6]), .Y(\MSG_TRP1_13_3_1_1[6] ));
    CFG4 #( .INIT(16'hFFFE) )  PRDATA30_2_0_sx_5 (.A(
        CoreAPB3_0_APBmslave3_PADDR[21]), .B(
        CoreAPB3_0_APBmslave3_PADDR[26]), .C(
        CoreAPB3_0_APBmslave3_PADDR[20]), .D(
        CoreAPB3_0_APBmslave3_PADDR[27]), .Y(PRDATA30_2_0_sx_5_net_1));
    SLE \MSG_WA_TRP1[4]  (.D(un1_PADDR_1_cry_4_S), .CLK(
        OSC_0_XTLOSC_O2F), .EN(N_986_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_MSG_WA_TRP1[4]));
    CFG4 #( .INIT(16'h0002) )  g2_5 (.A(
        CoreAPB3_0_APBmslave3_PADDR[29]), .B(
        CoreAPB3_0_APBmslave3_PADDR[7]), .C(
        CoreAPB3_0_APBmslave3_PADDR[13]), .D(
        CoreAPB3_0_APBmslave3_PADDR[0]), .Y(g2_5_net_1));
    SLE \APB_ADDRESS[31]  (.D(CoreAPB3_0_APBmslave3_PADDR[31]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[31]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  un25_TXB_0_o2_0 (.A(
        un25_TXB_0_o2_0_0_net_1), .B(un25_TXB_0_o2_0_1_net_1), .C(
        un25_TXB_0_o2_0_2_net_1), .D(un25_TXB_0_o2_0_3_net_1), .Y(
        N_982));
    CFG4 #( .INIT(16'h0001) )  PRDATA33_3 (.A(
        CoreAPB3_0_APBmslave3_PADDR[14]), .B(
        CoreAPB3_0_APBmslave3_PADDR[0]), .C(
        CoreAPB3_0_APBmslave3_PADDR[1]), .D(
        CoreAPB3_0_APBmslave3_PADDR[13]), .Y(PRDATA33_3_net_1));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[24]  (.A(
        COREEDAC_1_DATA_OUT[0]), .B(\PRDATA_14_0_iv_0_1[24]_net_1 ), 
        .C(un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[24] ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv[11]  (.A(
        COREEDAC_1_DATA_OUT[19]), .B(\PRDATA_14_0_iv_1[11]_net_1 ), .C(
        un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[11] ));
    CFG4 #( .INIT(16'hFFF2) )  Flag_Int_1_sqmuxa_1_i_0_0_1 (.A(
        pos1_Flag_A_HDL_Rec_Finish_net_1), .B(
        pos2_Flag_A_HDL_Rec_Finish_net_1), .C(
        Flag_Int_1_sqmuxa_1_i_0_0_1_0_net_1), .D(Flag_B_Rx18_net_1), 
        .Y(un1_Flag_Int_1_sqmuxa_1));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[10]  (.A(
        COREEDAC_1_DATA_OUT[18]), .B(\PRDATA_14_0_iv_0_sx[10]_net_1 ), 
        .C(\PRDATA_14_0_iv_0_1[10]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[10] ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv[20]  (.A(
        COREEDAC_1_DATA_OUT[12]), .B(\PRDATA_14_0_iv_1[20]_net_1 ), .C(
        un1_N_5_mux_0_0), .D(un1_N_5_mux_2), .Y(\PRDATA_14[20] ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_0_iv_0_0[14]  (.A(
        CLTU_0_TC_Packet_Counter[14]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(N_536), .Y(
        \PRDATA_14_0_iv_0_0[14]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  g0_3_4 (.A(
        CoreAPB3_0_APBmslave3_PADDR[11]), .B(
        CoreAPB3_0_APBmslave3_PADDR[7]), .C(
        CoreAPB3_0_APBmslave3_PADDR[12]), .D(
        CoreAPB3_0_APBmslave3_PADDR[13]), .Y(g0_3_4_net_1));
    SLE \MSG_TRP1[4]  (.D(\MSG_TRP1_13[4] ), .CLK(OSC_0_XTLOSC_O2F), 
        .EN(N_986_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(Glue_Logic_0_MSG_TRP1[4]));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[30]  (.A(
        COREEDAC_1_DATA_OUT[6]), .B(un1_N_5_mux_0_0), .C(
        \PRDATA_14_0_iv_0_1[30]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[30] ));
    SLE \PRDATA[28]  (.D(\PRDATA_14[28] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[28]));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_1[19]  (.A(PRDATA34_2_0)
        , .B(CLTU_0_TC_Error_Counter[19]), .C(
        \PRDATA_14_0_iv_1_1[19]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_1[19]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_0_iv_0_a3[30]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[30]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(N_563));
    CFG4 #( .INIT(16'h007F) )  PRDATA_N_5_mux_0_i_RNO (.A(
        CLTU_0_TC_Packet_Counter[4]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(N_618), .Y(PRDATA_m2_0_a2_2));
    SLE \MSG_WA_TRP1[7]  (.D(un1_PADDR_1_cry_7_S), .CLK(
        OSC_0_XTLOSC_O2F), .EN(N_986_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_MSG_WA_TRP1[7]));
    CFG4 #( .INIT(16'hFFFE) )  PRDATA30_2_0_sx_2 (.A(
        CoreAPB3_0_APBmslave3_PADDR[21]), .B(
        CoreAPB3_0_APBmslave3_PADDR[26]), .C(
        CoreAPB3_0_APBmslave3_PADDR[20]), .D(
        CoreAPB3_0_APBmslave3_PADDR[27]), .Y(PRDATA30_2_0_sx_2_net_1));
    CFG4 #( .INIT(16'hD5C0) )  \PRDATA_14_0_iv_0_sx_RNO[9]  (.A(N_982), 
        .B(PRDATA34_2_0), .C(un1_PRDATA30_4_0_a3_0_3), .D(
        Flag_m3_e_1_1), .Y(un1_PRDATA30_4_0_o3_sx));
    CFG4 #( .INIT(16'hFFFE) )  \APB_ADDRESS_RNILC92[10]  (.A(
        un1_PRDATA30_4_0_o3_0_11), .B(un1_PRDATA30_4_0_o3_0_14), .C(
        un1_PRDATA30_4_0_o3_0_13), .D(un1_PRDATA30_4_0_o3_0_12), .Y(
        N_1406));
    CFG4 #( .INIT(16'h0401) )  un1_PRDATA30_4_0_a3_0_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[2]), .B(
        CoreAPB3_0_APBmslave3_PADDR[4]), .C(
        CoreAPB3_0_APBmslave3_PADDR[5]), .D(
        CoreAPB3_0_APBmslave3_PADDR[3]), .Y(un1_PRDATA30_4_0_a3_0));
    CFG3 #( .INIT(8'h7F) )  un1_PRDATA47_1_i_0_o2_0 (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        CoreAPB3_0_APBmslave3_PENABLE), .C(iPSELS_raw23), .Y(N_977));
    CFG4 #( .INIT(16'h0015) )  PRDATA33_RNIO8525 (.A(N_651), .B(
        PRDATA34_2_0), .C(un1_PRDATA30_4_0_a3_0_3), .D(PRDATA33_net_1), 
        .Y(un1_m2_e_1));
    CFG4 #( .INIT(16'h195D) )  \MSG_TRP1_RNO_0[3]  (.A(
        \Byte_Count[1]_net_1 ), .B(\Byte_Count[0]_net_1 ), .C(
        CoreAPB3_0_APBmslave3_PWDATA[27]), .D(
        CoreAPB3_0_APBmslave3_PWDATA[11]), .Y(
        \MSG_TRP1_13_3_i_m2_1_1[3] ));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_iv_2_RNO[1]  (.A(
        CLTU_0_TC_Error_Counter[1]), .B(PRDATA34_2_0), .C(
        PRDATA38_1_0_net_1), .Y(\TC_Error_Counter_m[1] ));
    CFG4 #( .INIT(16'hF8FF) )  \PRDATA_14_iv_2[6]  (.A(PRDATA30), .B(
        CLTU_0_Flag_RX_ing), .C(\PRDATA_14_iv_0[6]_net_1 ), .D(
        \PRDATA_14_iv_2_1[6]_net_1 ), .Y(\PRDATA_14_iv_2[6]_net_1 ));
    SLE \PRDATA[16]  (.D(\PRDATA_14[16] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[16]));
    CFG4 #( .INIT(16'hFFFE) )  un25_TXB_0_o2_0_3 (.A(
        CoreAPB3_0_APBmslave3_PADDR[30]), .B(
        CoreAPB3_0_APBmslave3_PADDR[18]), .C(
        CoreAPB3_0_APBmslave3_PADDR[31]), .D(
        CoreAPB3_0_APBmslave3_PADDR[19]), .Y(un25_TXB_0_o2_0_3_net_1));
    CFG4 #( .INIT(16'h0020) )  un1_PRDATA30_4_0_o3_4_1_sx (.A(
        un1_PRDATA30_4_0_a3_0), .B(un1_PRDATA30_4_0_o3_4_sx_sx_0_net_1)
        , .C(PRDATA30_26_3), .D(un1_PRDATA30_4_0_o3_4_1_sx_sx_net_1), 
        .Y(un1_PRDATA30_4_0_o3_4_1_0));
    CFG3 #( .INIT(8'h39) )  \un1_APB_ADDRESS_3_1.SUM_i_x3[3]  (.A(
        un1_N_5_mux_2), .B(\APB_ADDRESS[5]_net_1 ), .C(N_644), .Y(
        N_49_i));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_0_1_1[28]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[28]), .B(
        CLTU_0_TC_Packet_Counter[28]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_0_1_1[28]_net_1 ));
    CFG4 #( .INIT(16'h0400) )  \PRDATA_14_iv_0_RNO_0[8]  (.A(
        CoreAPB3_0_APBmslave3_PADDR[2]), .B(
        CoreAPB3_0_APBmslave3_PADDR[4]), .C(
        CoreAPB3_0_APBmslave3_PADDR[5]), .D(
        CoreAPB3_0_APBmslave3_PADDR[3]), .Y(PRDATA_m1_0_a2_0));
    CFG4 #( .INIT(16'h8A00) )  \PRDATA_14_0_iv_0_sx[10]  (.A(
        PRDATA_m2_0), .B(N_660), .C(N_651), .D(N_629), .Y(
        \PRDATA_14_0_iv_0_sx[10]_net_1 ));
    SLE \PRDATA[21]  (.D(\PRDATA_14[21] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[21]));
    CFG3 #( .INIT(8'hBF) )  un1_PRDATA39_1_0_o3_1 (.A(
        \APB_ADDRESS[15]_net_1 ), .B(\APB_ADDRESS[14]_net_1 ), .C(
        \APB_ADDRESS[13]_net_1 ), .Y(N_644));
    SLE \PRDATA[22]  (.D(\PRDATA_14[22] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[22]));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv[13]  (.A(
        COREEDAC_1_DATA_OUT[21]), .B(\PRDATA_14_0_iv_1[13]_net_1 ), .C(
        un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[13] ));
    SLE \APB_ADDRESS[21]  (.D(CoreAPB3_0_APBmslave3_PADDR[21]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[21]_net_1 ));
    CFG4 #( .INIT(16'h0040) )  PRDATA36_2 (.A(
        CoreAPB3_0_APBmslave3_PADDR[1]), .B(
        CoreAPB3_0_APBmslave3_PADDR[29]), .C(
        CoreAPB3_0_APBmslave3_PADDR[28]), .D(
        CoreAPB3_0_APBmslave3_PADDR[0]), .Y(PRDATA36_2_net_1));
    CFG4 #( .INIT(16'hCCEC) )  Flag_B_Rx_0_sqmuxa_1_i_0_0 (.A(
        CoreAPB3_0_APBmslave3_PENABLE), .B(Flag_B_Rx18_net_1), .C(
        Flag_Int_0_sqmuxa_2_net_1), .D(CoreAPB3_0_APBmslave3_PWDATA[3])
        , .Y(Flag_B_Rx_0_sqmuxa_1_i_0_0_net_1));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_0_1[28]  (.A(
        PRDATA34_2_0), .B(CLTU_0_TC_Error_Counter[28]), .C(
        \PRDATA_14_0_iv_0_1_1[28]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_0_1[28]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un1_PADDR_1_cry_8 (.A(VCC_net_1), .B(
        CoreAPB3_0_APBmslave3_PADDR[8]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un1_PADDR_1_cry_7_net_1), .S(un1_PADDR_1_cry_8_S), .Y(), 
        .FCO(un1_PADDR_1_cry_8_net_1));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_14_iv_1_sx[0]  (.A(
        PRDATA30_2_0_4_net_1), .B(CLTU_0_TC_Error_Counter[0]), .C(
        PRDATA38_1_0_net_1), .D(PRDATA30_2_0_x_net_1), .Y(
        \PRDATA_14_iv_1_sx[0]_net_1 ));
    CFG4 #( .INIT(16'hFFF9) )  PRDATA33_1_0_0_o2_RNILO6E1 (.A(
        CoreAPB3_0_APBmslave3_PADDR[13]), .B(
        CoreAPB3_0_APBmslave3_PADDR[14]), .C(N_980), .D(N_982), .Y(
        N_984));
    SLE \APB_ADDRESS[27]  (.D(CoreAPB3_0_APBmslave3_PADDR[27]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[27]_net_1 ));
    CFG4 #( .INIT(16'h195D) )  \MSG_TRP1_RNO_0[1]  (.A(
        \Byte_Count[1]_net_1 ), .B(\Byte_Count[0]_net_1 ), .C(
        CoreAPB3_0_APBmslave3_PWDATA[25]), .D(
        CoreAPB3_0_APBmslave3_PWDATA[9]), .Y(
        \MSG_TRP1_13_3_i_m2_1_1[1] ));
    CFG3 #( .INIT(8'h80) )  Flag_Enable_1_sqmuxa_1_i_a2 (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        CoreAPB3_0_APBmslave3_PWRITE), .C(iPSELS_raw23), .Y(N_138));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[28]  (.A(
        COREEDAC_1_DATA_OUT[4]), .B(\PRDATA_14_0_iv_0_1[28]_net_1 ), 
        .C(un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[28] ));
    CFG4 #( .INIT(16'h80FF) )  \PRDATA_14_iv_0[3]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[3]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .D(\PRDATA_14_iv_0_1[3]_net_1 ), .Y(
        \PRDATA_14_iv_0[3]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \PRDATA_14_iv_0_o2_0_x_RNO[4]  (.A(
        CoreAPB3_0_APBmslave3_PADDR[7]), .B(
        CoreAPB3_0_APBmslave3_PADDR[11]), .C(
        CoreAPB3_0_APBmslave3_PADDR[13]), .Y(
        \PRDATA_14_iv_0_o2_0_x_RNO[4]_net_1 ));
    CFG3 #( .INIT(8'hAE) )  \PRDATA_14_0_iv_0_1[30]  (.A(
        \PRDATA_14_0_iv_0_0[30]_net_1 ), .B(
        CLTU_0_TC_Error_Counter[30]), .C(N_507), .Y(
        \PRDATA_14_0_iv_0_1[30]_net_1 ));
    CFG4 #( .INIT(16'h4657) )  \MSG_TRP1_RNO_0[0]  (.A(
        \Byte_Count[1]_net_1 ), .B(\Byte_Count[0]_net_1 ), .C(
        CoreAPB3_0_APBmslave3_PWDATA[16]), .D(
        CoreAPB3_0_APBmslave3_PWDATA[0]), .Y(
        \MSG_TRP1_13_3_i_m2_1_1[0] ));
    SLE \APB_ADDRESS[25]  (.D(CoreAPB3_0_APBmslave3_PADDR[25]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[25]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  un1_PRDATA30_4_0_o3_4_sx_sx_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[6]), .B(
        CoreAPB3_0_APBmslave3_PADDR[9]), .C(
        CoreAPB3_0_APBmslave3_PADDR[10]), .D(
        CoreAPB3_0_APBmslave3_PADDR[8]), .Y(
        un1_PRDATA30_4_0_o3_4_sx_sx_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_PADDR_1_cry_3 (.A(VCC_net_1), .B(
        CoreAPB3_0_APBmslave3_PADDR[3]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un1_PADDR_1_cry_2_net_1), .S(un1_PADDR_1_cry_3_S), .Y(), 
        .FCO(un1_PADDR_1_cry_3_net_1));
    ARI1 #( .INIT(20'h523DC) )  un1_PADDR_1_cry_1 (.A(
        CoreAPB3_0_APBmslave3_PADDR[1]), .B(\Byte_Count[0]_net_1 ), .C(
        \Byte_Count[1]_net_1 ), .D(N_984), .FCI(
        un1_PADDR_1_cry_0_net_1), .S(un1_PADDR_1_cry_1_S), .Y(), .FCO(
        un1_PADDR_1_cry_1_net_1));
    CFG3 #( .INIT(8'h04) )  \PRDATA_14_0_iv_0_sx_sx[9]  (.A(
        un1_m2_e_2_2_1_0), .B(N_651), .C(un1_PRDATA30_4_0_o3_4_0), .Y(
        \PRDATA_14_0_iv_0_sx_sx[9]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_iv_2_RNO[3]  (.A(
        CLTU_0_TC_Packet_Counter[3]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .Y(\TC_Packet_Counter_m[3] ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[26]  (.A(
        COREEDAC_1_DATA_OUT[2]), .B(\PRDATA_14_0_iv_0_1[26]_net_1 ), 
        .C(un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[26] ));
    CFG4 #( .INIT(16'h3B38) )  \MSG_TRP1_RNO[7]  (.A(
        CoreAPB3_0_APBmslave3_PWDATA[7]), .B(
        \MSG_TRP1_13_3_i_m2_1_1[7] ), .C(\Byte_Count[1]_net_1 ), .D(
        CoreAPB3_0_APBmslave3_PWDATA[15]), .Y(N_990));
    CFG4 #( .INIT(16'h8F88) )  \PRDATA_14_iv_0_sx[7]  (.A(
        un1_PRDATA30_4_0_a3_0_3), .B(PRDATA34_2_0), .C(
        un1_PRDATA30_4_0_o3_4), .D(un1_m2_e_2), .Y(
        \PRDATA_14_iv_0_sx[7]_net_1 ));
    CFG4 #( .INIT(16'hA8AA) )  PRDATA36_3_RNICLNN6 (.A(PRDATA34_2_0), 
        .B(PRDATA37_2_net_1), .C(PRDATA36_3_net_1), .D(
        un1_PRDATA30_4_0_o3_4_2), .Y(un1_PRDATA30_4_0_o3_4));
    SLE \MSG_WA_TRP1[0]  (.D(un1_PADDR_1_cry_0_Y), .CLK(
        OSC_0_XTLOSC_O2F), .EN(N_986_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_MSG_WA_TRP1[0]));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_iv_0_1_1_0[7]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[7]), .B(
        CLTU_0_TC_Packet_Counter[7]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_iv_0_1_1_0[7]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_iv_0_RNO[6]  (.A(
        CLTU_0_TC_Error_Counter[6]), .B(PRDATA34_2_0), .C(
        PRDATA38_1_0_net_1), .Y(\TC_Error_Counter_m[6] ));
    SLE \PRDATA[9]  (.D(\PRDATA_14[9] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[9]));
    SLE \APB_ADDRESS[14]  (.D(CoreAPB3_0_APBmslave3_PADDR[14]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[14]_net_1 ));
    CFG3 #( .INIT(8'hEA) )  \PRDATA_14_iv_0_2[7]  (.A(
        \PRDATA_14_iv_0_1[7] ), .B(Glue_Logic_0_Flag_Int_0[0]), .C(
        PRDATA30), .Y(\PRDATA_14_iv_0_2[7]_net_1 ));
    SLE \MSG_TRP1[2]  (.D(N_992), .CLK(OSC_0_XTLOSC_O2F), .EN(
        N_986_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(Glue_Logic_0_MSG_TRP1[2]));
    SLE \USER_RA_TRP1[2]  (.D(\APB_ADDRESS[4]_net_1 ), .CLK(
        OSC_0_XTLOSC_O2F), .EN(Flag_Enable_1_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_USER_RA_TRP1_1[2]));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_iv_0_RNO[1]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[1]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(\TM_Packet_Counter_m[1] ));
    GND GND (.Y(GND_net_1));
    SLE \APB_ADDRESS[10]  (.D(CoreAPB3_0_APBmslave3_PADDR[10]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[10]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_0_iv_0_a3[9]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[9]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(N_528));
    SLE \PRDATA[25]  (.D(\PRDATA_14[25] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[25]));
    CFG4 #( .INIT(16'hFFFE) )  un25_TXB_0_o2_0_2 (.A(
        CoreAPB3_0_APBmslave3_PADDR[21]), .B(
        CoreAPB3_0_APBmslave3_PADDR[26]), .C(
        CoreAPB3_0_APBmslave3_PADDR[20]), .D(
        CoreAPB3_0_APBmslave3_PADDR[27]), .Y(un25_TXB_0_o2_0_2_net_1));
    CFG4 #( .INIT(16'h0008) )  un1_PRDATA30_4_0_a3_0_4 (.A(
        un1_PRDATA30_4_0_a3_0_1), .B(PRDATA30_26_3), .C(
        un1_PRDATA30_4_0_a3_0_sx_0_net_1), .D(
        un1_PRDATA30_4_0_a3_0_4_sx_net_1), .Y(un1_PRDATA30_4_0_a3_0_3));
    CFG3 #( .INIT(8'h80) )  PRDATA30_2_0_x (.A(PRDATA30_2_0_2_net_1), 
        .B(PRDATA30_2_0_1_net_1), .C(PRDATA30_2_0_3_net_1), .Y(
        PRDATA30_2_0_x_net_1));
    CFG4 #( .INIT(16'h0100) )  Flag_Enable_RNIDIIB1 (.A(
        CoreAPB3_0_APBmslave3_PWRITE), .B(N_977), .C(Flag_Enable_net_1)
        , .D(N_651), .Y(Flag_Enable_RNIDIIB1_net_1));
    CFG4 #( .INIT(16'h0001) )  PRDATA30_2_0_2 (.A(
        CoreAPB3_0_APBmslave3_PADDR[23]), .B(
        CoreAPB3_0_APBmslave3_PADDR[24]), .C(
        CoreAPB3_0_APBmslave3_PADDR[25]), .D(
        CoreAPB3_0_APBmslave3_PADDR[22]), .Y(PRDATA30_2_0_2_net_1));
    CFG4 #( .INIT(16'h0004) )  PRDATA33 (.A(un25_TXB_0_o2_0_x_net_1), 
        .B(PRDATA33_6_net_1), .C(un25_TXB_0_o2_0_3_net_1), .D(N_980), 
        .Y(PRDATA33_net_1));
    SLE pos2_Flag_A_Tx_Finish (.D(pos1_Flag_A_Tx_Finish_net_1), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pos2_Flag_A_Tx_Finish_net_1));
    CFG4 #( .INIT(16'h4000) )  PRDATA33_6_x_RNI6QSC (.A(
        PRDATA33_1_0_0_o2_x_net_1), .B(Flag_m3_e_1_1_1), .C(
        PRDATA33_1_0_0_o2_1_net_1), .D(PRDATA33_4_net_1), .Y(
        Flag_m3_e_1_1));
    CFG4 #( .INIT(16'hFF04) )  Flag_Enable_1_sqmuxa_1_i_0 (.A(
        un1_PRDATA30_4_0_o3_4), .B(Flag_m1_e_1), .C(Flag_Enable_net_1), 
        .D(N_1000), .Y(Flag_Enable_1_sqmuxa_1_i_0_net_1));
    CFG4 #( .INIT(16'h8000) )  un1_PRDATA30_1_0_0_a2_0_a3 (.A(
        PRDATA34_26), .B(PRDATA34_2_0), .C(PRDATA30_1_0_0_a3_0_net_1), 
        .D(PRDATA35_1_0_0_a3_1_net_1), .Y(PRDATA30));
    SLE \MSG_WA_TRP1[3]  (.D(un1_PADDR_1_cry_3_S), .CLK(
        OSC_0_XTLOSC_O2F), .EN(N_986_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_MSG_WA_TRP1[3]));
    SLE \APB_ADDRESS[19]  (.D(CoreAPB3_0_APBmslave3_PADDR[19]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[19]_net_1 ));
    CFG4 #( .INIT(16'h7FFF) )  PRDATA38_1_0_0_RNI121D2 (.A(
        PRDATA37_1_0), .B(PRDATA30_26_4), .C(PRDATA38_1_0_0_net_1), .D(
        PRDATA30_26_3), .Y(g0_1_net_1));
    SLE \MSG_WA_TRP1[6]  (.D(un1_PADDR_1_cry_6_S), .CLK(
        OSC_0_XTLOSC_O2F), .EN(N_986_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_MSG_WA_TRP1[6]));
    CFG4 #( .INIT(16'h4450) )  PREADY_RNO_0 (.A(N_977), .B(
        PREADY_9_0_0_tz_net_1), .C(N_1025), .D(
        CoreAPB3_0_APBmslave3_PWRITE), .Y(un1_PRDATA47_1_i_0_a2_1_0));
    CFG4 #( .INIT(16'h5400) )  PRDATA_N_5_mux_0_i_1 (.A(PRDATA30), .B(
        N_660), .C(N_651), .D(PRDATA_m2_0_a2_0), .Y(
        PRDATA_N_5_mux_0_i_1_net_1));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv[15]  (.A(
        COREEDAC_1_DATA_OUT[23]), .B(un1_N_5_mux_0_0), .C(
        \PRDATA_14_0_iv_1[15]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[15] ));
    SLE \APB_ADDRESS[22]  (.D(CoreAPB3_0_APBmslave3_PADDR[22]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[22]_net_1 ));
    CFG3 #( .INIT(8'hEF) )  \PRDATA_14_iv_0_o2_0_x[4]  (.A(
        \PRDATA_14_iv_0_o2_0_0[4]_net_1 ), .B(
        CoreAPB3_0_APBmslave3_PADDR[12]), .C(
        \PRDATA_14_iv_0_o2_0_x_RNO[4]_net_1 ), .Y(
        \PRDATA_14_iv_0_o2_0_x[4]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  un25_TXB_0_o2_0_1 (.A(
        CoreAPB3_0_APBmslave3_PADDR[23]), .B(
        CoreAPB3_0_APBmslave3_PADDR[24]), .C(
        CoreAPB3_0_APBmslave3_PADDR[25]), .D(
        CoreAPB3_0_APBmslave3_PADDR[22]), .Y(un25_TXB_0_o2_0_1_net_1));
    CFG4 #( .INIT(16'hFFEC) )  \PRDATA_14_iv_2[2]  (.A(PRDATA30), .B(
        \PRDATA_14_iv_0[2]_net_1 ), .C(Flag_RX), .D(
        \TC_Error_Counter_m[2] ), .Y(\PRDATA_14_iv_2[2]_net_1 ));
    CFG4 #( .INIT(16'hFBFF) )  \PRDATA_14_iv_0_o2_0[4]  (.A(
        \PRDATA_14_iv_0_o2_0_0[4]_net_1 ), .B(PRDATA30_26_3), .C(
        \PRDATA_14_iv_0_o2_1_1[4]_net_1 ), .D(PRDATA30_26_4), .Y(N_510)
        );
    SLE \PRDATA[18]  (.D(\PRDATA_14[18] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[18]));
    SLE \APB_ADDRESS[23]  (.D(CoreAPB3_0_APBmslave3_PADDR[23]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[23]_net_1 ));
    CFG3 #( .INIT(8'hDC) )  PREADY_9_0_0_tz (.A(\Byte_Count[0]_net_1 ), 
        .B(N_984), .C(\Byte_Count[1]_net_1 ), .Y(PREADY_9_0_0_tz_net_1)
        );
    CFG4 #( .INIT(16'hFFFE) )  PRDATA30_2_0_sx_3 (.A(
        CoreAPB3_0_APBmslave3_PADDR[30]), .B(
        CoreAPB3_0_APBmslave3_PADDR[18]), .C(
        CoreAPB3_0_APBmslave3_PADDR[31]), .D(
        CoreAPB3_0_APBmslave3_PADDR[19]), .Y(PRDATA30_2_0_sx_3_net_1));
    SLE \USER_RA_TRP1[0]  (.D(\APB_ADDRESS[2]_net_1 ), .CLK(
        OSC_0_XTLOSC_O2F), .EN(Flag_Enable_1_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_USER_RA_TRP1_1[0]));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_1_1[19]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[19]), .B(
        CLTU_0_TC_Packet_Counter[19]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_1_1[19]_net_1 ));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_0_1[29]  (.A(
        PRDATA34_2_0), .B(CLTU_0_TC_Error_Counter[29]), .C(
        \PRDATA_14_0_iv_0_1_1[29]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_0_1[29]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  PRDATA38_i_o3 (.A(PRDATA38_1_0_net_1), .B(
        PRDATA30_2_0_4_net_1), .C(PRDATA30_2_0_x_net_1), .Y(N_507));
    CFG4 #( .INIT(16'h3B38) )  \MSG_TRP1_RNO[2]  (.A(
        CoreAPB3_0_APBmslave3_PWDATA[2]), .B(
        \MSG_TRP1_13_3_i_m2_1_1[2] ), .C(\Byte_Count[0]_net_1 ), .D(
        CoreAPB3_0_APBmslave3_PWDATA[18]), .Y(N_992));
    CFG3 #( .INIT(8'hAE) )  \PRDATA_14_0_iv_0_1[14]  (.A(
        \PRDATA_14_0_iv_0_0[14]_net_1 ), .B(
        CLTU_0_TC_Error_Counter[14]), .C(N_507), .Y(
        \PRDATA_14_0_iv_0_1[14]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_14_iv_0_2_sx[8]  (.A(
        PRDATA30_2_0_4_net_1), .B(CLTU_0_TC_Error_Counter[8]), .C(
        PRDATA38_1_0_net_1), .D(PRDATA30_2_0_x_net_1), .Y(
        \PRDATA_14_iv_0_2_sx[8]_net_1 ));
    SLE \APB_ADDRESS[5]  (.D(CoreAPB3_0_APBmslave3_PADDR[5]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[5]_net_1 ));
    SLE \APB_ADDRESS[26]  (.D(CoreAPB3_0_APBmslave3_PADDR[26]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[26]_net_1 ));
    SLE \PRDATA[7]  (.D(\PRDATA_14[7] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[7]));
    SLE \PRDATA[11]  (.D(\PRDATA_14[11] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[11]));
    CFG4 #( .INIT(16'hFEFA) )  \PRDATA_14_iv_2[1]  (.A(
        \TC_Error_Counter_m[1] ), .B(Glue_Logic_0_Flag_B_Tx), .C(
        \PRDATA_14_iv_0[1]_net_1 ), .D(PRDATA30), .Y(
        \PRDATA_14_iv_2[1]_net_1 ));
    SLE \PRDATA[12]  (.D(\PRDATA_14[12] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[12]));
    CFG4 #( .INIT(16'hAAA6) )  \Byte_Count_RNO[1]  (.A(
        \Byte_Count[1]_net_1 ), .B(\Byte_Count[0]_net_1 ), .C(N_985), 
        .D(N_984), .Y(N_1029_i_0));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_0_iv_0_a3_0[10]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[10]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(N_524));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv[22]  (.A(
        COREEDAC_1_DATA_OUT[14]), .B(\PRDATA_14_0_iv_1[22]_net_1 ), .C(
        un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[22] ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_0_iv_0_0[18]  (.A(
        CLTU_0_TC_Packet_Counter[18]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(N_540), .Y(
        \PRDATA_14_0_iv_0_0[18]_net_1 ));
    SLE \PRDATA[29]  (.D(\PRDATA_14[29] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[29]));
    SLE pos2_Flag_B_HDL_Rec_Finish (.D(
        pos1_Flag_B_HDL_Rec_Finish_net_1), .CLK(OSC_0_XTLOSC_O2F), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(pos2_Flag_B_HDL_Rec_Finish_net_1));
    CFG4 #( .INIT(16'hEFFF) )  PRDATA33_1_0_0_o2 (.A(
        CoreAPB3_0_APBmslave3_PADDR[10]), .B(
        CoreAPB3_0_APBmslave3_PADDR[12]), .C(PRDATA33_1_0_0_o2_1_net_1)
        , .D(CoreAPB3_0_APBmslave3_PADDR[28]), .Y(N_980));
    CFG4 #( .INIT(16'h80A0) )  \PRDATA_14_0_iv_0_sx[9]  (.A(N_629), .B(
        un1_PRDATA30_4_0_o3_sx), .C(PRDATA_m2_0), .D(
        \PRDATA_14_0_iv_0_sx_sx[9]_net_1 ), .Y(
        \PRDATA_14_0_iv_0_sx[9]_net_1 ));
    CFG4 #( .INIT(16'h4505) )  \PRDATA_14_iv_0_o2_0_RNIR1C82[4]  (.A(
        un1_PRDATA30_4_0_o3_4_0_sx), .B(un1_PRDATA30_4_0_a3_0), .C(
        N_510), .D(N_658), .Y(un1_PRDATA30_4_0_o3_4_0));
    SLE \PRDATA[6]  (.D(\PRDATA_14[6] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[6]));
    CFG4 #( .INIT(16'h0002) )  PRDATA30_2_0 (.A(PRDATA30_2_0_1_net_1), 
        .B(PRDATA30_2_0_sx_6_net_1), .C(PRDATA30_2_0_sx_4_net_1), .D(
        PRDATA30_2_0_sx_5_net_1), .Y(PRDATA34_2_0));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_iv_0_RNO[31]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[31]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(\TM_Packet_Counter_m[31] ));
    CFG4 #( .INIT(16'hFFAC) )  \PRDATA_14_iv_0[8]  (.A(
        COREEDAC_1_DATA_OUT[16]), .B(PRDATA_m1_0_a2_2), .C(
        un1_PRDATA39_1), .D(\PRDATA_14_iv_0_3[8]_net_1 ), .Y(
        \PRDATA_14[8] ));
    CFG4 #( .INIT(16'h3B38) )  \MSG_TRP1_RNO[3]  (.A(
        CoreAPB3_0_APBmslave3_PWDATA[3]), .B(
        \MSG_TRP1_13_3_i_m2_1_1[3] ), .C(\Byte_Count[0]_net_1 ), .D(
        CoreAPB3_0_APBmslave3_PWDATA[19]), .Y(N_991));
    SLE \PRDATA[24]  (.D(\PRDATA_14[24] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[24]));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_1[20]  (.A(PRDATA34_2_0)
        , .B(CLTU_0_TC_Error_Counter[20]), .C(
        \PRDATA_14_0_iv_1_1[20]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_1[20]_net_1 ));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_1[11]  (.A(PRDATA34_2_0)
        , .B(CLTU_0_TC_Error_Counter[11]), .C(
        \PRDATA_14_0_iv_1_1[11]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_1[11]_net_1 ));
    CFG3 #( .INIT(8'h20) )  PRDATA30_2_0_x_0 (.A(PRDATA30_2_0_2_net_1), 
        .B(PRDATA30_2_0_sx_0_net_1), .C(PRDATA30_2_0_1_net_1), .Y(
        PRDATA30_2_0_x_0_net_1));
    CFG4 #( .INIT(16'h8F0F) )  Flag_B_Tx_0_sqmuxa_1_i (.A(
        CoreAPB3_0_APBmslave3_PENABLE), .B(Flag_Int_0_sqmuxa_2_net_1), 
        .C(Flag_B_Tx18_net_1), .D(CoreAPB3_0_APBmslave3_PWDATA[1]), .Y(
        Flag_B_Tx_0_sqmuxa_1_i_0));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h0040) )  un25_TXB_0_o2_0_RNICK67D (.A(N_977), .B(
        N_651), .C(Flag_m3_e_1), .D(un1_m2_e_2_2_1_0), .Y(Flag_m1_e_1));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_iv[6]  (.A(
        COREEDAC_1_DATA_OUT[30]), .B(\PRDATA_14_iv_2[6]_net_1 ), .C(
        \PRDATA_14_iv_sx[6]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[6] ));
    CFG4 #( .INIT(16'hAA8A) )  PRDATA38_1_0_RNI2TOUI (.A(
        un1_PRDATA47_1_i_0_a2_0), .B(un1_PRDATA30_4_0_o3_0), .C(
        un1_PRDATA47_1_i_0_a2_1), .D(un1_PRDATA30_4_0_o3_4), .Y(
        un1_PRDATA47_1_i_0));
    SLE pos2_Flag_A_HDL_Rec_Finish (.D(
        pos1_Flag_A_HDL_Rec_Finish_net_1), .CLK(OSC_0_XTLOSC_O2F), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(pos2_Flag_A_HDL_Rec_Finish_net_1));
    CFG4 #( .INIT(16'h0001) )  g0_4 (.A(
        CoreAPB3_0_APBmslave3_PADDR[11]), .B(
        CoreAPB3_0_APBmslave3_PADDR[7]), .C(
        CoreAPB3_0_APBmslave3_PADDR[12]), .D(
        CoreAPB3_0_APBmslave3_PADDR[13]), .Y(PRDATA30_26_3));
    CFG4 #( .INIT(16'hEFFF) )  PRDATA30_2_0_x_0_RNIC2A05 (.A(
        PRDATA30_2_0_sx_net_1), .B(un1_PRDATA30_4_0_a3_0_4_sx_net_1), 
        .C(PRDATA30_2_0_x_0_net_1), .D(un1_PRDATA30_4_0_a3_0_4_x_net_1)
        , .Y(un1_m2_e_2_2_1));
    SLE \MSG_WA_TRP1[5]  (.D(un1_PADDR_1_cry_5_S), .CLK(
        OSC_0_XTLOSC_O2F), .EN(N_986_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_MSG_WA_TRP1[5]));
    CFG4 #( .INIT(16'hFFBF) )  un1_PRDATA30_4_0_o3_4_1_sx_sx (.A(
        CoreAPB3_0_APBmslave3_PADDR[1]), .B(
        CoreAPB3_0_APBmslave3_PADDR[29]), .C(
        CoreAPB3_0_APBmslave3_PADDR[28]), .D(
        CoreAPB3_0_APBmslave3_PADDR[0]), .Y(
        un1_PRDATA30_4_0_o3_4_1_sx_sx_net_1));
    CFG3 #( .INIT(8'hF4) )  \PRDATA_14_iv_1[0]  (.A(
        \PRDATA_14_iv_1_1[0]_net_1 ), .B(PRDATA34_2_0), .C(
        \PRDATA_14_iv_1_sx[0]_net_1 ), .Y(\PRDATA_14_iv_1[0]_net_1 ));
    SLE \PRDATA[15]  (.D(\PRDATA_14[15] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[15]));
    CFG3 #( .INIT(8'h15) )  PRDATA35_1_0_0_a3_RNIV4QV (.A(
        PRDATA38_1_0_net_1), .B(PRDATA30_1_0_0_a3_0_net_1), .C(N_658), 
        .Y(PRDATA35_1_0_0_a3_RNIV4QV_net_1));
    CFG4 #( .INIT(16'h0040) )  PRDATA36_1 (.A(
        CoreAPB3_0_APBmslave3_PADDR[2]), .B(
        CoreAPB3_0_APBmslave3_PADDR[4]), .C(
        CoreAPB3_0_APBmslave3_PADDR[5]), .D(
        CoreAPB3_0_APBmslave3_PADDR[3]), .Y(PRDATA36_1_net_1));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_0_iv_0_0[30]  (.A(
        CLTU_0_TC_Packet_Counter[30]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(N_563), .Y(
        \PRDATA_14_0_iv_0_0[30]_net_1 ));
    SLE Flag_B_Tx (.D(Flag_B_Tx18_net_1), .CLK(OSC_0_XTLOSC_O2F), .EN(
        Flag_B_Tx_0_sqmuxa_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_Flag_B_Tx));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_0_1_1[27]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[27]), .B(
        CLTU_0_TC_Packet_Counter[27]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_0_1_1[27]_net_1 ));
    CFG4 #( .INIT(16'hFFA2) )  PREADY_RNO (.A(un1_PRDATA47_1_i_0_a2_0), 
        .B(un1_m2_e_0_1), .C(un1_PRDATA30_4_0_o3_4), .D(
        un1_PRDATA47_1_i_0_a2_1_0), .Y(PREADY_9));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_1_1[11]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[11]), .B(
        CLTU_0_TC_Packet_Counter[11]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_1_1[11]_net_1 ));
    CFG4 #( .INIT(16'h8F0F) )  Flag_A_Tx_0_sqmuxa_1_i (.A(
        CoreAPB3_0_APBmslave3_PENABLE), .B(Flag_Int_0_sqmuxa_2_net_1), 
        .C(Flag_A_Tx18_net_1), .D(CoreAPB3_0_APBmslave3_PWDATA[0]), .Y(
        Flag_A_Tx_0_sqmuxa_1_i_0));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_0_1[21]  (.A(
        PRDATA34_2_0), .B(CLTU_0_TC_Error_Counter[21]), .C(
        \PRDATA_14_0_iv_0_1_1[21]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_0_1[21]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv[19]  (.A(
        COREEDAC_1_DATA_OUT[11]), .B(\PRDATA_14_0_iv_1[19]_net_1 ), .C(
        un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[19] ));
    CFG4 #( .INIT(16'h0200) )  Flag_Enable_RNI04AIK (.A(Flag_m3_e_1), 
        .B(un1_PRDATA30_4_0_o3_4), .C(un1_m2_e_2_2_1_0), .D(
        Flag_Enable_RNIDIIB1_net_1), .Y(Flag_Enable_1_sqmuxa));
    SLE \APB_ADDRESS[11]  (.D(CoreAPB3_0_APBmslave3_PADDR[11]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[11]_net_1 ));
    SLE \APB_ADDRESS[17]  (.D(CoreAPB3_0_APBmslave3_PADDR[17]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[17]_net_1 ));
    CFG4 #( .INIT(16'hD5C0) )  un25_TXB_0_o2_0_RNIO8SD5 (.A(N_982), .B(
        PRDATA34_2_0), .C(un1_PRDATA30_4_0_a3_0_3), .D(Flag_m3_e_1_1), 
        .Y(un1_PRDATA30_4_0_o3_0));
    ARI1 #( .INIT(20'h4AAA6) )  un1_PADDR_1_s_9 (.A(N_982), .B(
        CoreAPB3_0_APBmslave3_PADDR[9]), .C(un25_TXB_0_a2_0_net_1), .D(
        N_980), .FCI(un1_PADDR_1_cry_8_net_1), .S(un1_PADDR_1_s_9_S), 
        .Y(), .FCO());
    CFG4 #( .INIT(16'h8000) )  Flag_Int_0_sqmuxa_2 (.A(PRDATA34_2_0), 
        .B(N_138), .C(PRDATA30_1_0_0_a3_0_net_1), .D(N_658), .Y(
        Flag_Int_0_sqmuxa_2_net_1));
    CFG4 #( .INIT(16'h2A3F) )  un25_TXB_0_o2_0_RNIO8SD5_1 (.A(N_982), 
        .B(PRDATA34_2_0), .C(un1_PRDATA30_4_0_a3_0_3), .D(
        Flag_m3_e_1_1), .Y(Flag_m3_e_1));
    CFG4 #( .INIT(16'h0080) )  PRDATA37_1 (.A(
        CoreAPB3_0_APBmslave3_PADDR[5]), .B(
        CoreAPB3_0_APBmslave3_PADDR[29]), .C(
        CoreAPB3_0_APBmslave3_PADDR[28]), .D(
        CoreAPB3_0_APBmslave3_PADDR[0]), .Y(PRDATA37_1_0));
    SLE \MSG_WA_TRP1[1]  (.D(un1_PADDR_1_cry_1_S), .CLK(
        OSC_0_XTLOSC_O2F), .EN(N_986_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_MSG_WA_TRP1[1]));
    CFG4 #( .INIT(16'h8000) )  PRDATA38_1_0 (.A(PRDATA37_1_0), .B(
        PRDATA30_26_4), .C(PRDATA38_1_0_0_net_1), .D(PRDATA30_26_3), 
        .Y(PRDATA38_1_0_net_1));
    CFG4 #( .INIT(16'hFFEF) )  \APB_ADDRESS_RNI33P[16]  (.A(
        \APB_ADDRESS[16]_net_1 ), .B(un1_PRDATA30_4_0_o3_0_10), .C(
        \APB_ADDRESS[29]_net_1 ), .D(\APB_ADDRESS[17]_net_1 ), .Y(
        un1_PRDATA30_4_0_o3_0_14));
    CFG2 #( .INIT(4'h8) )  Flag_Enable1_RNIVHUL (.A(Flag_Enable_net_1), 
        .B(Flag_Enable1_net_1), .Y(N_1025));
    SLE \APB_ADDRESS[15]  (.D(CoreAPB3_0_APBmslave3_PADDR[15]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[15]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[29]  (.A(
        COREEDAC_1_DATA_OUT[5]), .B(\PRDATA_14_0_iv_0_1[29]_net_1 ), 
        .C(un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[29] ));
    CFG4 #( .INIT(16'hF4F0) )  Flag_Int_1_sqmuxa_1_i_0_0 (.A(
        CoreAPB3_0_APBmslave3_PWDATA[7]), .B(Flag_Int_0_sqmuxa_2_net_1)
        , .C(un1_Flag_Int_1_sqmuxa_1), .D(
        CoreAPB3_0_APBmslave3_PENABLE), .Y(
        Flag_Int_1_sqmuxa_1_i_0_0_net_1));
    CFG2 #( .INIT(4'h7) )  PRDATA30_2_0_RNIUQLC2 (.A(PRDATA34_2_0), .B(
        PRDATA34_26), .Y(PRDATA30_2_0_RNIUQLC2_net_1));
    SLE USER_REN_TRP1 (.D(Flag_Enable_i_0), .CLK(OSC_0_XTLOSC_O2F), 
        .EN(USER_REN_TRP1ce_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_USER_REN_TRP1));
    SLE \APB_ADDRESS[28]  (.D(CoreAPB3_0_APBmslave3_PADDR[28]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[28]_net_1 ));
    CFG2 #( .INIT(4'h4) )  PRDATA33_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[7]), .B(
        CoreAPB3_0_APBmslave3_PADDR[3]), .Y(PRDATA33_0_net_1));
    CFG4 #( .INIT(16'h193B) )  \MSG_TRP1_RNO_0[2]  (.A(
        \Byte_Count[0]_net_1 ), .B(\Byte_Count[1]_net_1 ), .C(
        CoreAPB3_0_APBmslave3_PWDATA[26]), .D(
        CoreAPB3_0_APBmslave3_PWDATA[10]), .Y(
        \MSG_TRP1_13_3_i_m2_1_1[2] ));
    CFG4 #( .INIT(16'hFFFE) )  \APB_ADDRESS_RNIQNG[24]  (.A(
        \APB_ADDRESS[27]_net_1 ), .B(\APB_ADDRESS[26]_net_1 ), .C(
        \APB_ADDRESS[25]_net_1 ), .D(\APB_ADDRESS[24]_net_1 ), .Y(
        un1_PRDATA30_4_0_o3_0_12));
    ARI1 #( .INIT(20'h4AA00) )  un1_PADDR_1_cry_2 (.A(VCC_net_1), .B(
        CoreAPB3_0_APBmslave3_PADDR[2]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un1_PADDR_1_cry_1_net_1), .S(un1_PADDR_1_cry_2_S), .Y(), 
        .FCO(un1_PADDR_1_cry_2_net_1));
    CFG4 #( .INIT(16'h0200) )  Flag_Enable1_1_sqmuxa_1_0_a2 (.A(
        Flag_Enable1_1_sqmuxa_1_1), .B(CoreAPB3_0_APBmslave3_PWRITE), 
        .C(un1_PRDATA30_4_0_o3_4), .D(Flag_m1_e_1), .Y(
        Flag_Enable1_1_sqmuxa_1));
    SLE \MSG_TRP1[7]  (.D(N_990), .CLK(OSC_0_XTLOSC_O2F), .EN(
        N_986_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(Glue_Logic_0_MSG_TRP1[7]));
    CFG4 #( .INIT(16'h1000) )  g0_3 (.A(CoreAPB3_0_APBmslave3_PADDR[9])
        , .B(CoreAPB3_0_APBmslave3_PADDR[6]), .C(g0_3_4_net_1), .D(
        g0_3_3_net_1), .Y(PRDATA34_26));
    CFG3 #( .INIT(8'h40) )  USER_REN_TRP1ce_1 (.A(
        CoreAPB3_0_APBmslave3_PWRITE), .B(
        CoreAPB3_0_APBmslave3_PENABLE), .C(iPSELS_raw23), .Y(
        USER_REN_TRP1ce_1_net_1));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_0_1[26]  (.A(
        PRDATA34_2_0), .B(CLTU_0_TC_Error_Counter[26]), .C(
        \PRDATA_14_0_iv_0_1_1[26]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_0_1[26]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_0_iv_0_a3[14]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[14]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(N_536));
    SLE \PRDATA[19]  (.D(\PRDATA_14[19] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[19]));
    SLE \MSG_TRP1[5]  (.D(\MSG_TRP1_13[5] ), .CLK(OSC_0_XTLOSC_O2F), 
        .EN(N_986_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(Glue_Logic_0_MSG_TRP1[5]));
    CFG4 #( .INIT(16'hFFBF) )  \PRDATA_14_iv_0_o2_1_1[4]  (.A(
        CoreAPB3_0_APBmslave3_PADDR[1]), .B(
        CoreAPB3_0_APBmslave3_PADDR[28]), .C(
        CoreAPB3_0_APBmslave3_PADDR[2]), .D(
        CoreAPB3_0_APBmslave3_PADDR[3]), .Y(
        \PRDATA_14_iv_0_o2_1_1[4]_net_1 ));
    CFG3 #( .INIT(8'hFB) )  PRDATA33_1_0_0_o2_x (.A(
        CoreAPB3_0_APBmslave3_PADDR[10]), .B(
        CoreAPB3_0_APBmslave3_PADDR[28]), .C(
        CoreAPB3_0_APBmslave3_PADDR[12]), .Y(PRDATA33_1_0_0_o2_x_net_1)
        );
    CFG2 #( .INIT(4'hD) )  Flag_A_Tx18 (.A(pos1_Flag_A_Tx_Finish_net_1)
        , .B(pos2_Flag_A_Tx_Finish_net_1), .Y(Flag_A_Tx18_net_1));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_0_1_1[26]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[26]), .B(
        CLTU_0_TC_Packet_Counter[26]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_0_1_1[26]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  PRDATA30_1_0_0_a3_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[2]), .B(
        CoreAPB3_0_APBmslave3_PADDR[4]), .C(
        CoreAPB3_0_APBmslave3_PADDR[5]), .D(
        CoreAPB3_0_APBmslave3_PADDR[3]), .Y(PRDATA30_1_0_0_a3_0_net_1));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv[23]  (.A(
        COREEDAC_1_DATA_OUT[15]), .B(un1_N_5_mux_0_0), .C(
        \PRDATA_14_0_iv_1[23]_net_1 ), .D(un1_N_5_mux_2), .Y(
        \PRDATA_14[23] ));
    CFG3 #( .INIT(8'h01) )  PRDATA33_3_x (.A(
        CoreAPB3_0_APBmslave3_PADDR[1]), .B(
        CoreAPB3_0_APBmslave3_PADDR[13]), .C(
        CoreAPB3_0_APBmslave3_PADDR[14]), .Y(PRDATA33_3_x_net_1));
    SLE \APB_ADDRESS[12]  (.D(CoreAPB3_0_APBmslave3_PADDR[12]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[12]_net_1 ));
    CFG4 #( .INIT(16'hFDFF) )  PRDATA30_2_0_sx_RNISNFN (.A(
        PRDATA30_2_0_2_net_1), .B(PRDATA30_2_0_sx_net_1), .C(
        PRDATA30_2_0_sx_0_net_1), .D(PRDATA30_2_0_1_net_1), .Y(
        un1_PRDATA30_4_0_o3_4_0_sx));
    SLE \PRDATA[14]  (.D(\PRDATA_14[14] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[14]));
    SLE \APB_ADDRESS[13]  (.D(CoreAPB3_0_APBmslave3_PADDR[13]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[13]_net_1 ));
    CFG4 #( .INIT(16'h0008) )  PRDATA37_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[4]), .B(
        CoreAPB3_0_APBmslave3_PADDR[2]), .C(
        CoreAPB3_0_APBmslave3_PADDR[3]), .D(
        CoreAPB3_0_APBmslave3_PADDR[1]), .Y(PRDATA37_0_net_1));
    CFG3 #( .INIT(8'hB3) )  PRDATA30_2_0_RNIVQVL4 (.A(
        un1_PRDATA30_4_0_a3_0_3), .B(N_651), .C(PRDATA34_2_0), .Y(
        un1_m2_e_0_1_sx));
    CFG3 #( .INIT(8'hAE) )  \PRDATA_14_0_iv_0_1[18]  (.A(
        \PRDATA_14_0_iv_0_0[18]_net_1 ), .B(
        CLTU_0_TC_Error_Counter[18]), .C(N_507), .Y(
        \PRDATA_14_0_iv_0_1[18]_net_1 ));
    CFG4 #( .INIT(16'h2F2C) )  \MSG_TRP1_RNO[5]  (.A(
        CoreAPB3_0_APBmslave3_PWDATA[5]), .B(\Byte_Count[1]_net_1 ), 
        .C(\MSG_TRP1_13_3_1_1[5] ), .D(
        CoreAPB3_0_APBmslave3_PWDATA[13]), .Y(\MSG_TRP1_13[5] ));
    CFG4 #( .INIT(16'hFFFD) )  \APB_ADDRESS_RNIC6D[10]  (.A(
        \APB_ADDRESS[28]_net_1 ), .B(\APB_ADDRESS[12]_net_1 ), .C(
        \APB_ADDRESS[11]_net_1 ), .D(\APB_ADDRESS[10]_net_1 ), .Y(
        un1_PRDATA30_4_0_o3_0_13));
    SLE Flag_Enable1 (.D(Flag_Enable1_1_sqmuxa_1), .CLK(
        OSC_0_XTLOSC_O2F), .EN(Flag_Enable1_1_sqmuxa_2_i_0_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Flag_Enable1_net_1));
    CFG4 #( .INIT(16'hFFFE) )  un1_PRDATA30_4_0_a3_0_sx_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[6]), .B(
        CoreAPB3_0_APBmslave3_PADDR[9]), .C(
        CoreAPB3_0_APBmslave3_PADDR[10]), .D(
        CoreAPB3_0_APBmslave3_PADDR[8]), .Y(
        un1_PRDATA30_4_0_a3_0_sx_0_net_1));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_0_1_1[24]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[24]), .B(
        CLTU_0_TC_Packet_Counter[24]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_0_1_1[24]_net_1 ));
    SLE \PRDATA[0]  (.D(\PRDATA_14[0] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[0]));
    CFG4 #( .INIT(16'hFF7F) )  PRDATA37_2_sx (.A(
        CoreAPB3_0_APBmslave3_PADDR[5]), .B(
        CoreAPB3_0_APBmslave3_PADDR[29]), .C(
        CoreAPB3_0_APBmslave3_PADDR[28]), .D(
        CoreAPB3_0_APBmslave3_PADDR[0]), .Y(PRDATA37_2_sx_net_1));
    CFG3 #( .INIT(8'h02) )  \PRDATA_14_iv_0_3_RNO[8]  (.A(
        un1_m2_e_2_2_1), .B(N_651), .C(PRDATA33_net_1), .Y(
        \PRDATA_14_iv_0_3_RNO[8]_net_1 ));
    SLE \PRDATA[31]  (.D(\PRDATA_14[31] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[31]));
    CFG1 #( .INIT(2'h1) )  USER_REN_TRP1_RNO (.A(Flag_Enable_net_1), 
        .Y(Flag_Enable_i_0));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_iv_0_RNO[2]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[2]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(\TM_Packet_Counter_m[2] ));
    SLE \APB_ADDRESS[16]  (.D(CoreAPB3_0_APBmslave3_PADDR[16]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[16]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  un25_TXB_0_o2_0_RNI8U09J (.A(
        un1_m2_e_2_2_1_0), .B(N_1406), .C(un1_PRDATA30_4_0_o3_4), .D(
        un1_PRDATA30_4_0_o3_0), .Y(un1_N_5_mux_2));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_1[12]  (.A(PRDATA34_2_0)
        , .B(CLTU_0_TC_Error_Counter[12]), .C(
        \PRDATA_14_0_iv_1_1[12]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_1[12]_net_1 ));
    CFG3 #( .INIT(8'hAE) )  \PRDATA_14_0_iv_1[15]  (.A(
        \PRDATA_14_0_iv_0[15]_net_1 ), .B(CLTU_0_TC_Error_Counter[15]), 
        .C(N_507), .Y(\PRDATA_14_0_iv_1[15]_net_1 ));
    SLE pos2_Flag_B_Tx_Finish (.D(pos1_Flag_B_Tx_Finish_net_1), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pos2_Flag_B_Tx_Finish_net_1));
    SLE \PRDATA[4]  (.D(PRDATA_N_5_mux_0_i_0), .CLK(OSC_0_XTLOSC_O2F), 
        .EN(un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[4]));
    CFG4 #( .INIT(16'hFFFE) )  PRDATA30_2_0_sx_4 (.A(
        CoreAPB3_0_APBmslave3_PADDR[23]), .B(
        CoreAPB3_0_APBmslave3_PADDR[24]), .C(
        CoreAPB3_0_APBmslave3_PADDR[25]), .D(
        CoreAPB3_0_APBmslave3_PADDR[22]), .Y(PRDATA30_2_0_sx_4_net_1));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_1_1[20]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[20]), .B(
        CLTU_0_TC_Packet_Counter[20]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_1_1[20]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_0_iv_0_RNO[23]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[23]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(\TM_Packet_Counter_m[23] ));
    CFG4 #( .INIT(16'hFF40) )  Flag_Enable1_1_sqmuxa_2_i_0 (.A(
        un1_PRDATA30_4_0_o3_4), .B(Flag_m1_e_1), .C(
        Flag_Enable1_1_sqmuxa_1_1), .D(N_1000), .Y(
        Flag_Enable1_1_sqmuxa_2_i_0_net_1));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_iv_1_1[0]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[0]), .B(
        CLTU_0_TC_Packet_Counter[0]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_iv_1_1[0]_net_1 ));
    CFG4 #( .INIT(16'h7FFF) )  PRDATA30_2_0_3_RNIUOJ6 (.A(
        PRDATA30_2_0_1_net_1), .B(PRDATA30_2_0_3_net_1), .C(
        PRDATA30_2_0_2_net_1), .D(PRDATA30_2_0_4_net_1), .Y(
        PRDATA30_2_0_3_RNIUOJ6_net_1));
    CFG4 #( .INIT(16'h337F) )  PRDATA_N_5_mux_0_i_1_RNO (.A(
        CLTU_0_TC_Error_Counter[4]), .B(PRDATA34_2_0), .C(
        PRDATA38_1_0_net_1), .D(un1_PRDATA30_4_0_a3_0_3), .Y(
        PRDATA_m2_0_a2_0));
    CFG4 #( .INIT(16'h0800) )  PRDATA37_2 (.A(PRDATA37_0_net_1), .B(
        PRDATA30_26_3), .C(PRDATA37_2_sx_net_1), .D(PRDATA30_26_4), .Y(
        PRDATA37_2_net_1));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_0_iv_0_0[9]  (.A(
        CLTU_0_TC_Packet_Counter[9]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(N_528), .Y(\PRDATA_14_0_iv_0_0[9]_net_1 )
        );
    CFG4 #( .INIT(16'h8F83) )  \MSG_TRP1_RNO[4]  (.A(
        CoreAPB3_0_APBmslave3_PWDATA[12]), .B(\Byte_Count[0]_net_1 ), 
        .C(\MSG_TRP1_13_3_1_1[4] ), .D(
        CoreAPB3_0_APBmslave3_PWDATA[28]), .Y(\MSG_TRP1_13[4] ));
    CFG3 #( .INIT(8'hFE) )  un25_TXB_0_o2_0_x (.A(
        un25_TXB_0_o2_0_0_net_1), .B(un25_TXB_0_o2_0_1_net_1), .C(
        un25_TXB_0_o2_0_2_net_1), .Y(un25_TXB_0_o2_0_x_net_1));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_1[13]  (.A(PRDATA34_2_0)
        , .B(CLTU_0_TC_Error_Counter[13]), .C(
        \PRDATA_14_0_iv_1_1[13]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_1[13]_net_1 ));
    SLE \PRDATA[20]  (.D(\PRDATA_14[20] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[20]));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_0_iv_0[15]  (.A(
        CLTU_0_TC_Packet_Counter[15]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(\TM_Packet_Counter_m[15] ), .Y(
        \PRDATA_14_0_iv_0[15]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  PRDATA33_RNIDN5GC (.A(un1_m2_e_2_2_1), 
        .B(un1_m2_e_2_2_1_0), .C(N_651), .D(PRDATA33_net_1), .Y(
        un1_m2_e_2));
    SLE \Byte_Count[1]  (.D(N_1029_i_0), .CLK(OSC_0_XTLOSC_O2F), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Byte_Count[1]_net_1 ));
    CFG4 #( .INIT(16'h8F88) )  \PRDATA_14_iv_sx[5]  (.A(
        un1_PRDATA30_4_0_a3_0_3), .B(PRDATA34_2_0), .C(
        un1_PRDATA30_4_0_o3_4), .D(un1_m2_e_2), .Y(
        \PRDATA_14_iv_sx[5]_net_1 ));
    SLE \PRDATA[2]  (.D(\PRDATA_14[2] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[2]));
    CFG4 #( .INIT(16'h0001) )  PRDATA33_4 (.A(
        CoreAPB3_0_APBmslave3_PADDR[5]), .B(
        CoreAPB3_0_APBmslave3_PADDR[4]), .C(
        CoreAPB3_0_APBmslave3_PADDR[6]), .D(
        CoreAPB3_0_APBmslave3_PADDR[9]), .Y(PRDATA33_4_net_1));
    CFG4 #( .INIT(16'h0001) )  PRDATA30_2_0_1 (.A(
        CoreAPB3_0_APBmslave3_PADDR[14]), .B(
        CoreAPB3_0_APBmslave3_PADDR[17]), .C(
        CoreAPB3_0_APBmslave3_PADDR[15]), .D(
        CoreAPB3_0_APBmslave3_PADDR[16]), .Y(PRDATA30_2_0_1_net_1));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv[25]  (.A(
        COREEDAC_1_DATA_OUT[1]), .B(\PRDATA_14_0_iv_1[25]_net_1 ), .C(
        un1_N_5_mux_0_0), .D(un1_N_5_mux_2), .Y(\PRDATA_14[25] ));
    SLE \MSG_WA_TRP1[9]  (.D(un1_PADDR_1_s_9_S), .CLK(OSC_0_XTLOSC_O2F)
        , .EN(N_986_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_MSG_WA_TRP1[9]));
    CFG4 #( .INIT(16'h00FB) )  \PRDATA_14_iv_0_o2_0_x_RNIQHN76[4]  (.A(
        \PRDATA_14_iv_0_o2_1_1[4]_net_1 ), .B(PRDATA30_26_4), .C(
        \PRDATA_14_iv_0_o2_0_x[4]_net_1 ), .D(
        un1_PRDATA30_4_0_o3_4_1_0), .Y(un1_PRDATA30_4_0_o3_4_2));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_0_1_1[21]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[21]), .B(
        CLTU_0_TC_Packet_Counter[21]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_0_1_1[21]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  USER_REN_TRP1ce (.A(un1_m2_e_0_1), .B(
        un1_PRDATA30_4_0_o3_4), .C(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .D(
        USER_REN_TRP1ce_1_net_1), .Y(USER_REN_TRP1ce_net_1));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_0_1_1[29]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[29]), .B(
        CLTU_0_TC_Packet_Counter[29]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_0_1_1[29]_net_1 ));
    CFG3 #( .INIT(8'hAE) )  \PRDATA_14_0_iv_1[17]  (.A(
        \PRDATA_14_0_iv_0[17]_net_1 ), .B(CLTU_0_TC_Error_Counter[17]), 
        .C(N_507), .Y(\PRDATA_14_0_iv_1[17]_net_1 ));
    CFG4 #( .INIT(16'h2F2C) )  \MSG_TRP1_RNO[1]  (.A(
        CoreAPB3_0_APBmslave3_PWDATA[1]), .B(\Byte_Count[0]_net_1 ), 
        .C(\MSG_TRP1_13_3_i_m2_1_1[1] ), .D(
        CoreAPB3_0_APBmslave3_PWDATA[17]), .Y(N_993));
    SLE \MSG_TRP1[1]  (.D(N_993), .CLK(OSC_0_XTLOSC_O2F), .EN(
        N_986_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(Glue_Logic_0_MSG_TRP1[1]));
    ARI1 #( .INIT(20'h4AA00) )  un1_PADDR_1_cry_4 (.A(VCC_net_1), .B(
        CoreAPB3_0_APBmslave3_PADDR[4]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un1_PADDR_1_cry_3_net_1), .S(un1_PADDR_1_cry_4_S), .Y(), 
        .FCO(un1_PADDR_1_cry_4_net_1));
    SLE Flag_A_Tx (.D(Flag_A_Tx18_net_1), .CLK(OSC_0_XTLOSC_O2F), .EN(
        Flag_A_Tx_0_sqmuxa_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        TXD4_net_0));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_0_iv_0_RNO[15]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[15]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(\TM_Packet_Counter_m[15] ));
    CFG3 #( .INIT(8'hFE) )  un25_TXB_0_o2_0_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[15]), .B(
        CoreAPB3_0_APBmslave3_PADDR[16]), .C(
        CoreAPB3_0_APBmslave3_PADDR[17]), .Y(un25_TXB_0_o2_0_0_net_1));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_iv_0_2_0[8]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[8]), .B(
        CLTU_0_TC_Packet_Counter[8]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_iv_0_2_0[8]_net_1 ));
    SLE \PRDATA[23]  (.D(\PRDATA_14[23] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[23]));
    CFG2 #( .INIT(4'h2) )  un25_TXB_0_a2_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[14]), .B(
        CoreAPB3_0_APBmslave3_PADDR[13]), .Y(un25_TXB_0_a2_0_net_1));
    SLE \PRDATA[8]  (.D(\PRDATA_14[8] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[8]));
    CFG4 #( .INIT(16'h193B) )  \MSG_TRP1_RNO_0[7]  (.A(
        \Byte_Count[1]_net_1 ), .B(\Byte_Count[0]_net_1 ), .C(
        CoreAPB3_0_APBmslave3_PWDATA[31]), .D(
        CoreAPB3_0_APBmslave3_PWDATA[23]), .Y(
        \MSG_TRP1_13_3_i_m2_1_1[7] ));
    SLE \APB_ADDRESS[3]  (.D(CoreAPB3_0_APBmslave3_PADDR[3]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[3]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_iv_0[2]  (.A(
        CLTU_0_TC_Packet_Counter[2]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(\TM_Packet_Counter_m[2] ), .Y(
        \PRDATA_14_iv_0[2]_net_1 ));
    SLE pos1_Flag_A_Tx_Finish (.D(CPU_W_HDL_R_0_Flag_A_Tx_Finish), 
        .CLK(OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pos1_Flag_A_Tx_Finish_net_1));
    CFG4 #( .INIT(16'h0001) )  g2_6 (.A(
        CoreAPB3_0_APBmslave3_PADDR[12]), .B(
        CoreAPB3_0_APBmslave3_PADDR[11]), .C(
        CoreAPB3_0_APBmslave3_PADDR[6]), .D(
        CoreAPB3_0_APBmslave3_PADDR[9]), .Y(g2_6_net_1));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_iv[0]  (.A(
        COREEDAC_1_DATA_OUT[24]), .B(un1_N_5_mux_0_0), .C(
        \PRDATA_14_iv_2[0]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[0] ));
    CFG4 #( .INIT(16'hFFFE) )  \APB_ADDRESS_RNICBI[22]  (.A(
        \APB_ADDRESS[31]_net_1 ), .B(\APB_ADDRESS[30]_net_1 ), .C(
        \APB_ADDRESS[23]_net_1 ), .D(\APB_ADDRESS[22]_net_1 ), .Y(
        un1_PRDATA30_4_0_o3_0_11));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_iv[5]  (.A(
        COREEDAC_1_DATA_OUT[29]), .B(\PRDATA_14_iv_2[5]_net_1 ), .C(
        \PRDATA_14_iv_sx[5]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[5] ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_0_iv_0[17]  (.A(
        CLTU_0_TC_Packet_Counter[17]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(\TM_Packet_Counter_m[17] ), .Y(
        \PRDATA_14_0_iv_0[17]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \APB_ADDRESS_RNIKFE[18]  (.A(
        \APB_ADDRESS[21]_net_1 ), .B(\APB_ADDRESS[20]_net_1 ), .C(
        \APB_ADDRESS[19]_net_1 ), .D(\APB_ADDRESS[18]_net_1 ), .Y(
        un1_PRDATA30_4_0_o3_0_10));
    CFG4 #( .INIT(16'hFFFD) )  \PRDATA_14_iv_0_o2_0_0[4]  (.A(
        CoreAPB3_0_APBmslave3_PADDR[29]), .B(
        CoreAPB3_0_APBmslave3_PADDR[4]), .C(
        CoreAPB3_0_APBmslave3_PADDR[5]), .D(
        CoreAPB3_0_APBmslave3_PADDR[0]), .Y(
        \PRDATA_14_iv_0_o2_0_0[4]_net_1 ));
    CFG3 #( .INIT(8'hC9) )  \Byte_Count_RNO[0]  (.A(N_984), .B(
        \Byte_Count[0]_net_1 ), .C(N_985), .Y(N_145_i_0));
    CFG4 #( .INIT(16'h1011) )  un25_TXB_0_o2_0_RNI0GIHC (.A(
        un1_m2_e_0_1_sx), .B(un1_m2_e_2_2_1_0), .C(N_982), .D(
        Flag_m3_e_1_1), .Y(un1_m2_e_0_1));
    CFG3 #( .INIT(8'h20) )  un1_PRDATA30_4_0_a3_0_4_x (.A(
        PRDATA30_26_3), .B(un1_PRDATA30_4_0_a3_0_sx_0_net_1), .C(
        un1_PRDATA30_4_0_a3_0_1), .Y(un1_PRDATA30_4_0_a3_0_4_x_net_1));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_iv[31]  (.A(
        COREEDAC_1_DATA_OUT[7]), .B(un1_N_5_mux_0_0), .C(
        \PRDATA_14_iv_2[31]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[31] ));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_0_iv_0_RNO[17]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[17]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(\TM_Packet_Counter_m[17] ));
    CFG4 #( .INIT(16'hFAFE) )  \PRDATA_14_iv_2[31]  (.A(PRDATA30), .B(
        CLTU_0_TC_Error_Counter[31]), .C(\PRDATA_14_iv_0[31]_net_1 ), 
        .D(N_507), .Y(\PRDATA_14_iv_2[31]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[21]  (.A(
        COREEDAC_1_DATA_OUT[13]), .B(\PRDATA_14_0_iv_0_1[21]_net_1 ), 
        .C(un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[21] ));
    CFG4 #( .INIT(16'h8F88) )  \PRDATA_14_iv_sx[3]  (.A(
        un1_PRDATA30_4_0_a3_0_3), .B(PRDATA34_2_0), .C(
        un1_PRDATA30_4_0_o3_4), .D(un1_m2_e_2), .Y(
        \PRDATA_14_iv_sx[3]_net_1 ));
    CFG4 #( .INIT(16'hCCEC) )  Flag_A_Rx_0_sqmuxa_1_i_0_0 (.A(
        CoreAPB3_0_APBmslave3_PENABLE), .B(Flag_A_Rx18_net_1), .C(
        Flag_Int_0_sqmuxa_2_net_1), .D(CoreAPB3_0_APBmslave3_PWDATA[2])
        , .Y(Flag_A_Rx_0_sqmuxa_1_i_0_0_net_1));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_0_iv_0_0[10]  (.A(
        CLTU_0_TC_Packet_Counter[10]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(N_524), .Y(
        \PRDATA_14_0_iv_0_0[10]_net_1 ));
    SLE \APB_ADDRESS[18]  (.D(CoreAPB3_0_APBmslave3_PADDR[18]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[18]_net_1 ));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_1_1[13]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[13]), .B(
        CLTU_0_TC_Packet_Counter[13]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_1_1[13]_net_1 ));
    SLE PREADY (.D(PREADY_9), .CLK(OSC_0_XTLOSC_O2F), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PREADY));
    CFG4 #( .INIT(16'hBF3F) )  PRDATA_N_5_mux_0_i (.A(
        COREEDAC_1_DATA_OUT[28]), .B(PRDATA_m2_0_a2_2), .C(
        PRDATA_N_5_mux_0_i_1_net_1), .D(un1_PRDATA39_1), .Y(
        PRDATA_N_5_mux_0_i_0));
    CFG4 #( .INIT(16'h7FFF) )  \PRDATA_14_iv_0_1[3]  (.A(
        PRDATA30_2_0_4_net_1), .B(CLTU_0_TC_Error_Counter[3]), .C(
        PRDATA38_1_0_net_1), .D(PRDATA30_2_0_x_net_1), .Y(
        \PRDATA_14_iv_0_1[3]_net_1 ));
    SLE pos1_Flag_B_HDL_Rec_Finish (.D(
        HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pos1_Flag_B_HDL_Rec_Finish_net_1));
    CFG4 #( .INIT(16'h193B) )  \MSG_TRP1_RNO_0[5]  (.A(
        \Byte_Count[1]_net_1 ), .B(\Byte_Count[0]_net_1 ), .C(
        CoreAPB3_0_APBmslave3_PWDATA[29]), .D(
        CoreAPB3_0_APBmslave3_PWDATA[21]), .Y(\MSG_TRP1_13_3_1_1[5] ));
    CFG3 #( .INIT(8'h7F) )  \PRDATA_14_iv_2_1[5]  (.A(
        CLTU_0_TC_Packet_Counter[5]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .Y(\PRDATA_14_iv_2_1[5]_net_1 ));
    SLE \Byte_Count[0]  (.D(N_145_i_0), .CLK(OSC_0_XTLOSC_O2F), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Byte_Count[0]_net_1 ));
    SLE \PRDATA[27]  (.D(\PRDATA_14[27] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[27]));
    SLE \PRDATA[1]  (.D(\PRDATA_14[1] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[1]));
    SLE \APB_ADDRESS[2]  (.D(CoreAPB3_0_APBmslave3_PADDR[2]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[2]_net_1 ));
    SLE \PRDATA[3]  (.D(\PRDATA_14[3] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[3]));
    CFG3 #( .INIT(8'h7F) )  \PRDATA_14_iv_2_1[6]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[6]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(\PRDATA_14_iv_2_1[6]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[9]  (.A(
        COREEDAC_1_DATA_OUT[17]), .B(\PRDATA_14_0_iv_0_sx[9]_net_1 ), 
        .C(\PRDATA_14_0_iv_0_1[9]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[9] ));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_0_1[27]  (.A(
        PRDATA34_2_0), .B(CLTU_0_TC_Error_Counter[27]), .C(
        \PRDATA_14_0_iv_0_1_1[27]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_0_1[27]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[14]  (.A(
        COREEDAC_1_DATA_OUT[22]), .B(un1_N_5_mux_0_0), .C(
        \PRDATA_14_0_iv_0_1[14]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[14] ));
    CFG4 #( .INIT(16'h0001) )  PRDATA30_2_0_3 (.A(
        CoreAPB3_0_APBmslave3_PADDR[21]), .B(
        CoreAPB3_0_APBmslave3_PADDR[26]), .C(
        CoreAPB3_0_APBmslave3_PADDR[20]), .D(
        CoreAPB3_0_APBmslave3_PADDR[27]), .Y(PRDATA30_2_0_3_net_1));
    SLE Flag_B_Rx (.D(Flag_B_Rx18_net_1), .CLK(OSC_0_XTLOSC_O2F), .EN(
        Flag_B_Rx_0_sqmuxa_1_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_Flag_B_Rx));
    CFG3 #( .INIT(8'hAE) )  \PRDATA_14_0_iv_0_1[9]  (.A(
        \PRDATA_14_0_iv_0_0[9]_net_1 ), .B(CLTU_0_TC_Error_Counter[9]), 
        .C(N_507), .Y(\PRDATA_14_0_iv_0_1[9]_net_1 ));
    CFG4 #( .INIT(16'h8F83) )  \MSG_TRP1_RNO[0]  (.A(
        CoreAPB3_0_APBmslave3_PWDATA[8]), .B(\Byte_Count[0]_net_1 ), 
        .C(\MSG_TRP1_13_3_i_m2_1_1[0] ), .D(
        CoreAPB3_0_APBmslave3_PWDATA[24]), .Y(N_994));
    SLE \MSG_TRP1[3]  (.D(N_991), .CLK(OSC_0_XTLOSC_O2F), .EN(
        N_986_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(Glue_Logic_0_MSG_TRP1[3]));
    CFG4 #( .INIT(16'h0210) )  \APB_ADDRESS_RNI3P7M[13]  (.A(
        \APB_ADDRESS[13]_net_1 ), .B(N_1025), .C(
        \APB_ADDRESS[15]_net_1 ), .D(\APB_ADDRESS[14]_net_1 ), .Y(
        \APB_ADDRESS_RNI3P7M[13]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  PRDATA30_2_0_4 (.A(
        CoreAPB3_0_APBmslave3_PADDR[30]), .B(
        CoreAPB3_0_APBmslave3_PADDR[18]), .C(
        CoreAPB3_0_APBmslave3_PADDR[31]), .D(
        CoreAPB3_0_APBmslave3_PADDR[19]), .Y(PRDATA30_2_0_4_net_1));
    SLE pos1_Flag_A_HDL_Rec_Finish (.D(
        HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        pos1_Flag_A_HDL_Rec_Finish_net_1));
    CFG4 #( .INIT(16'h4000) )  PRDATA33_6 (.A(
        CoreAPB3_0_APBmslave3_PADDR[8]), .B(PRDATA33_0_net_1), .C(
        PRDATA33_3_net_1), .D(PRDATA33_4_net_1), .Y(PRDATA33_6_net_1));
    SLE \PRDATA[10]  (.D(\PRDATA_14[10] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[10]));
    CFG4 #( .INIT(16'h0020) )  PRDATA38_1_0_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[4]), .B(
        CoreAPB3_0_APBmslave3_PADDR[2]), .C(
        CoreAPB3_0_APBmslave3_PADDR[3]), .D(
        CoreAPB3_0_APBmslave3_PADDR[1]), .Y(PRDATA38_1_0_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un1_PADDR_1_cry_6 (.A(VCC_net_1), .B(
        CoreAPB3_0_APBmslave3_PADDR[6]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un1_PADDR_1_cry_5_net_1), .S(un1_PADDR_1_cry_6_S), .Y(), 
        .FCO(un1_PADDR_1_cry_6_net_1));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_iv_2_RNO[2]  (.A(
        CLTU_0_TC_Error_Counter[2]), .B(PRDATA34_2_0), .C(
        PRDATA38_1_0_net_1), .Y(\TC_Error_Counter_m[2] ));
    CFG4 #( .INIT(16'h0001) )  g0_5 (.A(CoreAPB3_0_APBmslave3_PADDR[6])
        , .B(CoreAPB3_0_APBmslave3_PADDR[9]), .C(
        CoreAPB3_0_APBmslave3_PADDR[10]), .D(
        CoreAPB3_0_APBmslave3_PADDR[8]), .Y(PRDATA30_26_4));
    SLE \MSG_TRP1[0]  (.D(N_994), .CLK(OSC_0_XTLOSC_O2F), .EN(
        N_986_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(Glue_Logic_0_MSG_TRP1[0]));
    CFG4 #( .INIT(16'h020F) )  PRDATA38_1_0_0_RNIFJ317 (.A(g2_8_net_1), 
        .B(N_506), .C(g0_sx), .D(g0_1_net_1), .Y(un1_m2_e_2_2_1_0));
    CFG4 #( .INIT(16'h8F83) )  \MSG_TRP1_RNO[6]  (.A(
        CoreAPB3_0_APBmslave3_PWDATA[14]), .B(\Byte_Count[0]_net_1 ), 
        .C(\MSG_TRP1_13_3_1_1[6] ), .D(
        CoreAPB3_0_APBmslave3_PWDATA[30]), .Y(\MSG_TRP1_13[6] ));
    CFG3 #( .INIT(8'hEA) )  \PRDATA_14_iv_2[0]  (.A(
        \PRDATA_14_iv_1[0]_net_1 ), .B(TXD4_net_0), .C(PRDATA30), .Y(
        \PRDATA_14_iv_2[0]_net_1 ));
    CFG4 #( .INIT(16'hFF7F) )  g0_1 (.A(
        CoreAPB3_0_APBmslave3_PADDR[28]), .B(
        CoreAPB3_0_APBmslave3_PADDR[3]), .C(PRDATA32_4), .D(
        g0_1_0_net_1), .Y(N_506));
    CFG2 #( .INIT(4'hD) )  Flag_B_Tx18 (.A(pos1_Flag_B_Tx_Finish_net_1)
        , .B(pos2_Flag_B_Tx_Finish_net_1), .Y(Flag_B_Tx18_net_1));
    CFG4 #( .INIT(16'hFFFE) )  PRDATA30_2_0_sx (.A(
        CoreAPB3_0_APBmslave3_PADDR[30]), .B(
        CoreAPB3_0_APBmslave3_PADDR[18]), .C(
        CoreAPB3_0_APBmslave3_PADDR[31]), .D(
        CoreAPB3_0_APBmslave3_PADDR[19]), .Y(PRDATA30_2_0_sx_net_1));
    CFG4 #( .INIT(16'h0004) )  un25_TXB_0_o2_0_RNIC5A9J (.A(
        un1_m2_e_2_2_1_0), .B(N_651), .C(un1_PRDATA30_4_0_o3_4), .D(
        un1_PRDATA30_4_0_o3_0), .Y(un1_PRDATA39_1));
    CFG2 #( .INIT(4'hE) )  g0_1_0 (.A(CoreAPB3_0_APBmslave3_PADDR[1]), 
        .B(CoreAPB3_0_APBmslave3_PADDR[2]), .Y(g0_1_0_net_1));
    CFG4 #( .INIT(16'h7FFF) )  PREADY_9_0_o2 (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        CoreAPB3_0_APBmslave3_PWRITE), .C(
        CoreAPB3_0_APBmslave3_PENABLE), .D(iPSELS_raw23), .Y(N_985));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_1_1[25]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[25]), .B(
        CLTU_0_TC_Packet_Counter[25]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_1_1[25]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv[17]  (.A(
        COREEDAC_1_DATA_OUT[9]), .B(un1_N_5_mux_0_0), .C(
        \PRDATA_14_0_iv_1[17]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[17] ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_iv[3]  (.A(
        COREEDAC_1_DATA_OUT[27]), .B(\PRDATA_14_iv_2[3]_net_1 ), .C(
        \PRDATA_14_iv_sx[3]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[3] ));
    CFG4 #( .INIT(16'h0210) )  \APB_ADDRESS_RNIPJI2[13]  (.A(
        \APB_ADDRESS[13]_net_1 ), .B(N_1406), .C(
        \APB_ADDRESS[15]_net_1 ), .D(\APB_ADDRESS[14]_net_1 ), .Y(
        N_651));
    ARI1 #( .INIT(20'h4AA00) )  un1_PADDR_1_cry_7 (.A(VCC_net_1), .B(
        CoreAPB3_0_APBmslave3_PADDR[7]), .C(GND_net_1), .D(GND_net_1), 
        .FCI(un1_PADDR_1_cry_6_net_1), .S(un1_PADDR_1_cry_7_S), .Y(), 
        .FCO(un1_PADDR_1_cry_7_net_1));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_iv_0[5]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[5]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .D(\TC_Error_Counter_m[5] ), .Y(
        \PRDATA_14_iv_0[5]_net_1 ));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_1_1[12]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[12]), .B(
        CLTU_0_TC_Packet_Counter[12]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_1_1[12]_net_1 ));
    SLE \PRDATA[13]  (.D(\PRDATA_14[13] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[13]));
    CFG4 #( .INIT(16'hFFF7) )  un1_PRDATA30_4_0_i_a2 (.A(PRDATA30_26_4)
        , .B(PRDATA30_26_3), .C(un1_PRDATA30_4_0_i_a2_1_0_net_1), .D(
        un1_PRDATA30_4_0_i_a2_sx_net_1), .Y(N_629));
    CFG4 #( .INIT(16'hF0F2) )  \PRDATA_14_iv_0_3[8]  (.A(
        \PRDATA_14_iv_0_3_RNO[8]_net_1 ), .B(un1_m2_e_2_2_1_0), .C(
        \PRDATA_14_iv_0_2[8]_net_1 ), .D(un1_PRDATA30_4_0_o3_4), .Y(
        \PRDATA_14_iv_0_3[8]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_0_iv_0_a3[18]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[18]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(N_540));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_0_1_1[16]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[16]), .B(
        CLTU_0_TC_Packet_Counter[16]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_0_1_1[16]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[18]  (.A(
        COREEDAC_1_DATA_OUT[10]), .B(un1_N_5_mux_0_0), .C(
        \PRDATA_14_0_iv_0_1[18]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[18] ));
    CFG4 #( .INIT(16'h1000) )  g2_8 (.A(CoreAPB3_0_APBmslave3_PADDR[8])
        , .B(CoreAPB3_0_APBmslave3_PADDR[10]), .C(g2_5_net_1), .D(
        g2_6_net_1), .Y(g2_8_net_1));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_iv_0_RNO[5]  (.A(
        CLTU_0_TC_Error_Counter[5]), .B(PRDATA34_2_0), .C(
        PRDATA38_1_0_net_1), .Y(\TC_Error_Counter_m[5] ));
    CFG4 #( .INIT(16'h135F) )  un1_PRDATA30_4_0_i_a2_1_0 (.A(
        PRDATA36_1_net_1), .B(PRDATA37_0_net_1), .C(PRDATA36_2_net_1), 
        .D(PRDATA37_1_0), .Y(un1_PRDATA30_4_0_i_a2_1_0_net_1));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_iv_0[1]  (.A(
        CLTU_0_TC_Packet_Counter[1]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(\TM_Packet_Counter_m[1] ), .Y(
        \PRDATA_14_iv_0[1]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  PRDATA30_2_0_sx_6 (.A(
        CoreAPB3_0_APBmslave3_PADDR[30]), .B(
        CoreAPB3_0_APBmslave3_PADDR[18]), .C(
        CoreAPB3_0_APBmslave3_PADDR[31]), .D(
        CoreAPB3_0_APBmslave3_PADDR[19]), .Y(PRDATA30_2_0_sx_6_net_1));
    SLE Flag_A_Rx (.D(Flag_A_Rx18_net_1), .CLK(OSC_0_XTLOSC_O2F), .EN(
        Flag_A_Rx_0_sqmuxa_1_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(Flag_RX));
    SLE \APB_ADDRESS[30]  (.D(CoreAPB3_0_APBmslave3_PADDR[30]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[30]_net_1 ));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_0_1[16]  (.A(
        PRDATA34_2_0), .B(CLTU_0_TC_Error_Counter[16]), .C(
        \PRDATA_14_0_iv_0_1_1[16]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_0_1[16]_net_1 ));
    CFG2 #( .INIT(4'h2) )  Flag_Enable1_1_sqmuxa_1_0_a2_1 (.A(
        Flag_Enable_net_1), .B(Flag_Enable1_net_1), .Y(
        Flag_Enable1_1_sqmuxa_1_1));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[16]  (.A(
        COREEDAC_1_DATA_OUT[8]), .B(\PRDATA_14_0_iv_0_1[16]_net_1 ), 
        .C(un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[16] ));
    SLE \MSG_TRP1[6]  (.D(\MSG_TRP1_13[6] ), .CLK(OSC_0_XTLOSC_O2F), 
        .EN(N_986_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(Glue_Logic_0_MSG_TRP1[6]));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_14_iv_0_RNO[8]  (.A(
        PRDATA_m1_0_a2_0), .B(PRDATA35_1_0_0_a3_1_net_1), .C(
        PRDATA34_26), .D(PRDATA34_2_0), .Y(PRDATA_m1_0_a2_2));
    CFG4 #( .INIT(16'hFFBF) )  un1_PRDATA30_4_0_a3_0_4_sx (.A(
        CoreAPB3_0_APBmslave3_PADDR[1]), .B(
        CoreAPB3_0_APBmslave3_PADDR[29]), .C(
        CoreAPB3_0_APBmslave3_PADDR[28]), .D(
        CoreAPB3_0_APBmslave3_PADDR[0]), .Y(
        un1_PRDATA30_4_0_a3_0_4_sx_net_1));
    CFG4 #( .INIT(16'hFEEE) )  \PRDATA_14_iv_2[3]  (.A(
        \TC_Packet_Counter_m[3] ), .B(\PRDATA_14_iv_0[3]_net_1 ), .C(
        Glue_Logic_0_Flag_B_Rx), .D(PRDATA30), .Y(
        \PRDATA_14_iv_2[3]_net_1 ));
    CFG3 #( .INIT(8'h80) )  \PRDATA_14_iv_0_a3_1[4]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[4]), .B(PRDATA34_2_0), .C(
        PRDATA36_3_net_1), .Y(N_618));
    CFG4 #( .INIT(16'h153F) )  \PRDATA_14_0_iv_1_1[22]  (.A(
        CPU_W_HDL_R_0_TM_Packet_Counter[22]), .B(
        CLTU_0_TC_Packet_Counter[22]), .C(PRDATA37_2_net_1), .D(
        PRDATA36_3_net_1), .Y(\PRDATA_14_0_iv_1_1[22]_net_1 ));
    CFG4 #( .INIT(16'h7FFF) )  PRDATA30_2_0_3_RNIUOJ6_0 (.A(
        PRDATA30_2_0_1_net_1), .B(PRDATA30_2_0_3_net_1), .C(
        PRDATA30_2_0_2_net_1), .D(PRDATA30_2_0_4_net_1), .Y(g0_sx));
    SLE \USER_RA_TRP1[3]  (.D(N_49_i), .CLK(OSC_0_XTLOSC_O2F), .EN(
        Flag_Enable_1_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_USER_RA_TRP1_1[3]));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_1[22]  (.A(PRDATA34_2_0)
        , .B(CLTU_0_TC_Error_Counter[22]), .C(
        \PRDATA_14_0_iv_1_1[22]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_1[22]_net_1 ));
    CFG2 #( .INIT(4'h2) )  Flag_A_Rx18 (.A(
        pos1_Flag_A_HDL_Rec_Finish_net_1), .B(
        pos2_Flag_A_HDL_Rec_Finish_net_1), .Y(Flag_A_Rx18_net_1));
    SLE \MSG_WA_TRP1[2]  (.D(un1_PADDR_1_cry_2_S), .CLK(
        OSC_0_XTLOSC_O2F), .EN(N_986_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_MSG_WA_TRP1[2]));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_1[25]  (.A(PRDATA34_2_0)
        , .B(CLTU_0_TC_Error_Counter[25]), .C(
        \PRDATA_14_0_iv_1_1[25]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_1[25]_net_1 ));
    CFG4 #( .INIT(16'h0A0E) )  PRDATA33_RNIUMP46 (.A(
        PRDATA30_2_0_RNIUQLC2_net_1), .B(
        PRDATA35_1_0_0_a3_RNIV4QV_net_1), .C(PRDATA33_net_1), .D(
        \PRDATA_14_iv_0_o2_1_RNI894C2[4]_net_1 ), .Y(PRDATA_m2_0));
    CFG4 #( .INIT(16'hFBFF) )  un1_PRDATA30_4_0_i_a2_sx (.A(
        PRDATA30_2_0_sx_2_net_1), .B(PRDATA30_2_0_1_net_1), .C(
        PRDATA30_2_0_sx_3_net_1), .D(PRDATA30_2_0_2_net_1), .Y(
        un1_PRDATA30_4_0_i_a2_sx_net_1));
    CFG4 #( .INIT(16'h0ACE) )  \PRDATA_14_0_iv_0_1[24]  (.A(
        PRDATA34_2_0), .B(CLTU_0_TC_Error_Counter[24]), .C(
        \PRDATA_14_0_iv_0_1_1[24]_net_1 ), .D(N_507), .Y(
        \PRDATA_14_0_iv_0_1[24]_net_1 ));
    CFG4 #( .INIT(16'h0203) )  PRDATA38_1_0_RNI1TLQ5 (.A(
        PRDATA30_2_0_3_RNIUOJ6_net_1), .B(N_1406), .C(
        un1_PRDATA47_1_i_0_a2_N_3L3_1), .D(PRDATA38_1_0_net_1), .Y(
        un1_PRDATA47_1_i_0_a2_1));
    CFG4 #( .INIT(16'hFFEF) )  un1_PRDATA30_4_0_i_a2_RNI73S6F (.A(
        un1_m2_e_2_2_1_0), .B(un1_PRDATA30_4_0_o3_sx_0), .C(N_629), .D(
        un1_PRDATA30_4_0_o3_4_0), .Y(N_660));
    CFG2 #( .INIT(4'h4) )  PRDATA33_1_0_0_o2_1 (.A(
        CoreAPB3_0_APBmslave3_PADDR[11]), .B(
        CoreAPB3_0_APBmslave3_PADDR[29]), .Y(PRDATA33_1_0_0_o2_1_net_1)
        );
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_iv[2]  (.A(
        COREEDAC_1_DATA_OUT[26]), .B(un1_N_5_mux_0_0), .C(
        \PRDATA_14_iv_2[2]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[2] ));
    SLE \PRDATA[17]  (.D(\PRDATA_14[17] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[17]));
    CFG4 #( .INIT(16'h5575) )  \APB_ADDRESS_RNIHAAA5[13]  (.A(
        \APB_ADDRESS_RNI3P7M[13]_net_1 ), .B(N_506), .C(g2_8_net_1), 
        .D(PRDATA30_2_0_3_RNIUOJ6_net_1), .Y(
        un1_PRDATA47_1_i_0_a2_N_3L3_1));
    CFG4 #( .INIT(16'h0040) )  PRDATA35_1_0_0_a3_1 (.A(
        CoreAPB3_0_APBmslave3_PADDR[1]), .B(
        CoreAPB3_0_APBmslave3_PADDR[29]), .C(
        CoreAPB3_0_APBmslave3_PADDR[28]), .D(
        CoreAPB3_0_APBmslave3_PADDR[0]), .Y(PRDATA35_1_0_0_a3_1_net_1));
    CFG4 #( .INIT(16'hD5C0) )  un25_TXB_0_o2_0_RNIO8SD5_0 (.A(N_982), 
        .B(PRDATA34_2_0), .C(un1_PRDATA30_4_0_a3_0_3), .D(
        Flag_m3_e_1_1), .Y(un1_PRDATA30_4_0_o3_sx_0));
    CFG4 #( .INIT(16'h8F88) )  \PRDATA_14_iv_sx[6]  (.A(
        un1_PRDATA30_4_0_a3_0_3), .B(PRDATA34_2_0), .C(
        un1_PRDATA30_4_0_o3_4), .D(un1_m2_e_2), .Y(
        \PRDATA_14_iv_sx[6]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv[12]  (.A(
        COREEDAC_1_DATA_OUT[20]), .B(\PRDATA_14_0_iv_1[12]_net_1 ), .C(
        un1_N_5_mux_0_0), .D(un1_N_5_mux_2), .Y(\PRDATA_14[12] ));
    SLE \APB_ADDRESS[4]  (.D(CoreAPB3_0_APBmslave3_PADDR[4]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[4]_net_1 ));
    CFG4 #( .INIT(16'h0040) )  un1_PRDATA30_4_0_i_a2_RNI735RE (.A(
        un1_m2_e_2_2_1_0), .B(un1_m2_e_1), .C(N_629), .D(
        un1_PRDATA30_4_0_o3_4_0), .Y(un1_N_5_mux_0_0));
    CFG3 #( .INIT(8'hAE) )  \PRDATA_14_0_iv_1[23]  (.A(
        \PRDATA_14_0_iv_0[23]_net_1 ), .B(CLTU_0_TC_Error_Counter[23]), 
        .C(N_507), .Y(\PRDATA_14_0_iv_1[23]_net_1 ));
    SLE \APB_ADDRESS[24]  (.D(CoreAPB3_0_APBmslave3_PADDR[24]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[24]_net_1 ));
    SLE USER_WEN_TRP1 (.D(VCC_net_1), .CLK(OSC_0_XTLOSC_O2F), .EN(
        N_986_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(Glue_Logic_0_USER_WEN_TRP1));
    CFG3 #( .INIT(8'hAE) )  \PRDATA_14_0_iv_0_1[10]  (.A(
        \PRDATA_14_0_iv_0_0[10]_net_1 ), .B(
        CLTU_0_TC_Error_Counter[10]), .C(N_507), .Y(
        \PRDATA_14_0_iv_0_1[10]_net_1 ));
    SLE \APB_ADDRESS[20]  (.D(CoreAPB3_0_APBmslave3_PADDR[20]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[20]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_iv_0[6]  (.A(
        CLTU_0_TC_Packet_Counter[6]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(\TC_Error_Counter_m[6] ), .Y(
        \PRDATA_14_iv_0[6]_net_1 ));
    ARI1 #( .INIT(20'h545BA) )  un1_PADDR_1_cry_0 (.A(
        CoreAPB3_0_APBmslave3_PADDR[0]), .B(\Byte_Count[0]_net_1 ), .C(
        \Byte_Count[1]_net_1 ), .D(N_984), .FCI(GND_net_1), .S(), .Y(
        un1_PADDR_1_cry_0_Y), .FCO(un1_PADDR_1_cry_0_net_1));
    SLE \PRDATA[26]  (.D(\PRDATA_14[26] ), .CLK(OSC_0_XTLOSC_O2F), .EN(
        un1_PRDATA47_1_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[26]));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_iv[1]  (.A(
        COREEDAC_1_DATA_OUT[25]), .B(un1_N_5_mux_0_0), .C(
        \PRDATA_14_iv_2[1]_net_1 ), .D(un1_PRDATA39_1), .Y(
        \PRDATA_14[1] ));
    CFG4 #( .INIT(16'h1000) )  PRDATA33_6_x (.A(
        CoreAPB3_0_APBmslave3_PADDR[0]), .B(
        CoreAPB3_0_APBmslave3_PADDR[8]), .C(PRDATA33_0_net_1), .D(
        PRDATA33_3_x_net_1), .Y(Flag_m3_e_1_1_1));
    CFG4 #( .INIT(16'h0008) )  un1_PRDATA30_4_0_a3_0_2 (.A(
        CoreAPB3_0_APBmslave3_PADDR[2]), .B(
        CoreAPB3_0_APBmslave3_PADDR[4]), .C(
        CoreAPB3_0_APBmslave3_PADDR[5]), .D(
        CoreAPB3_0_APBmslave3_PADDR[3]), .Y(un1_PRDATA30_4_0_a3_0_1));
    CFG2 #( .INIT(4'hB) )  \PRDATA_14_iv_0_o2_1[4]  (.A(
        \PRDATA_14_iv_0_o2_1_1[4]_net_1 ), .B(PRDATA32_4), .Y(N_502));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_0_iv_0[23]  (.A(
        CLTU_0_TC_Packet_Counter[23]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(\TM_Packet_Counter_m[23] ), .Y(
        \PRDATA_14_0_iv_0[23]_net_1 ));
    CFG4 #( .INIT(16'hECCC) )  Flag_Enable_1_sqmuxa_1_i_o2 (.A(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        CoreAPB3_0_APBmslave3_PREADY), .C(iPSELS_raw23), .D(
        CoreAPB3_0_APBmslave3_PWRITE), .Y(N_1000));
    CFG4 #( .INIT(16'h0222) )  \PRDATA_14_iv_0_o2_1_RNI894C2[4]  (.A(
        CoreAPB3_0_APBmslave3_PADDR[29]), .B(
        CoreAPB3_0_APBmslave3_PADDR[0]), .C(N_506), .D(N_502), .Y(
        \PRDATA_14_iv_0_o2_1_RNI894C2[4]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_14_iv_0[31]  (.A(
        CLTU_0_TC_Packet_Counter[31]), .B(PRDATA34_2_0), .C(
        PRDATA37_2_net_1), .D(\TM_Packet_Counter_m[31] ), .Y(
        \PRDATA_14_iv_0[31]_net_1 ));
    CFG4 #( .INIT(16'h2637) )  \MSG_TRP1_RNO_0[4]  (.A(
        \Byte_Count[0]_net_1 ), .B(\Byte_Count[1]_net_1 ), .C(
        CoreAPB3_0_APBmslave3_PWDATA[20]), .D(
        CoreAPB3_0_APBmslave3_PWDATA[4]), .Y(\MSG_TRP1_13_3_1_1[4] ));
    CFG3 #( .INIT(8'h80) )  PRDATA35_1_0_0_a3 (.A(PRDATA30_26_4), .B(
        PRDATA30_26_3), .C(PRDATA35_1_0_0_a3_1_net_1), .Y(N_658));
    CFG2 #( .INIT(4'h1) )  g0_3_3 (.A(CoreAPB3_0_APBmslave3_PADDR[10]), 
        .B(CoreAPB3_0_APBmslave3_PADDR[8]), .Y(g0_3_3_net_1));
    CFG2 #( .INIT(4'h1) )  g0_2 (.A(CoreAPB3_0_APBmslave3_PADDR[5]), 
        .B(CoreAPB3_0_APBmslave3_PADDR[4]), .Y(PRDATA32_4));
    SLE \APB_ADDRESS[29]  (.D(CoreAPB3_0_APBmslave3_PADDR[29]), .CLK(
        OSC_0_XTLOSC_O2F), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \APB_ADDRESS[29]_net_1 ));
    CFG2 #( .INIT(4'h2) )  Flag_B_Rx18 (.A(
        pos1_Flag_B_HDL_Rec_Finish_net_1), .B(
        pos2_Flag_B_HDL_Rec_Finish_net_1), .Y(Flag_B_Rx18_net_1));
    SLE \Flag_Int_1[0]  (.D(un1_Flag_Int_1_sqmuxa_1), .CLK(
        OSC_0_XTLOSC_O2F), .EN(Flag_Int_1_sqmuxa_1_i_0_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Glue_Logic_0_Flag_Int_0[0]));
    CFG4 #( .INIT(16'hBFAA) )  \PRDATA_14_iv_0_2[8]  (.A(
        \PRDATA_14_iv_0_2_sx[8]_net_1 ), .B(
        \PRDATA_14_iv_0_2_0[8]_net_1 ), .C(N_510), .D(PRDATA34_2_0), 
        .Y(\PRDATA_14_iv_0_2[8]_net_1 ));
    CFG4 #( .INIT(16'hFEFC) )  \PRDATA_14_0_iv_0[27]  (.A(
        COREEDAC_1_DATA_OUT[3]), .B(\PRDATA_14_0_iv_0_1[27]_net_1 ), 
        .C(un1_N_5_mux_0_0), .D(un1_PRDATA39_1), .Y(\PRDATA_14[27] ));
    
endmodule


module Convolutional_Encoder(
       shift1_reg_4,
       shift1_reg_0,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       P_CLK,
       c_in,
       Convolutional_Encoder_out_1_0
    );
output shift1_reg_4;
output shift1_reg_0;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  P_CLK;
input  c_in;
output Convolutional_Encoder_out_1_0;

    wire \shift1_reg[5]_net_1 , VCC_net_1, GND_net_1, 
        \shift1_reg[3]_net_1 , \shift1_reg[2]_net_1 , 
        \shift1_reg[1]_net_1 ;
    
    SLE \shift1_reg[4]  (.D(\shift1_reg[3]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(shift1_reg_4));
    SLE \shift1_reg[0]  (.D(c_in), .CLK(P_CLK), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        shift1_reg_0));
    VCC VCC (.Y(VCC_net_1));
    SLE \shift1_reg[3]  (.D(\shift1_reg[2]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\shift1_reg[3]_net_1 ));
    SLE \shift1_reg[5]  (.D(shift1_reg_4), .CLK(P_CLK), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \shift1_reg[5]_net_1 ));
    SLE \shift1_reg[2]  (.D(\shift1_reg[1]_net_1 ), .CLK(P_CLK), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\shift1_reg[2]_net_1 ));
    SLE \shift1_reg[1]  (.D(shift1_reg_0), .CLK(P_CLK), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \shift1_reg[1]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  Convolutional_Encoder_out_0_0 (.A(c_in), 
        .B(\shift1_reg[5]_net_1 ), .C(\shift1_reg[2]_net_1 ), .D(
        \shift1_reg[1]_net_1 ), .Y(Convolutional_Encoder_out_1_0));
    
endmodule


module test_4463andcpuopration_COREEDAC_0_actram(
       CODE_FROM_RAM,
       Bit_Count_16dec_i_1,
       CODED,
       Glue_Logic_0_MSG_TRP1,
       Glue_Logic_0_MSG_WA_TRP1,
       CPU_W_HDL_R_0_USER_RA_TRP1_0,
       CPU_W_HDL_R_0_USER_RA_TRP1_1,
       CPU_W_HDL_R_0_USER_RA_TRP1_2,
       CPU_W_HDL_R_0_USER_RA_TRP1_3,
       CPU_W_HDL_R_0_USER_RA_TRP1_4,
       CPU_W_HDL_R_0_USER_RA_TRP1_5,
       CPU_W_HDL_R_0_USER_RA_TRP1_6,
       CPU_W_HDL_R_0_USER_RA_TRP1_7,
       CPU_W_HDL_R_0_USER_RA_TRP1_9,
       CPU_W_HDL_R_0_USER_REN_TRP1,
       OSC_0_XTLOSC_O2F,
       Glue_Logic_0_USER_WEN_TRP1
    );
output [12:0] CODE_FROM_RAM;
input  [3:3] Bit_Count_16dec_i_1;
input  [4:0] CODED;
input  [7:0] Glue_Logic_0_MSG_TRP1;
input  [9:0] Glue_Logic_0_MSG_WA_TRP1;
input  CPU_W_HDL_R_0_USER_RA_TRP1_0;
input  CPU_W_HDL_R_0_USER_RA_TRP1_1;
input  CPU_W_HDL_R_0_USER_RA_TRP1_2;
input  CPU_W_HDL_R_0_USER_RA_TRP1_3;
input  CPU_W_HDL_R_0_USER_RA_TRP1_4;
input  CPU_W_HDL_R_0_USER_RA_TRP1_5;
input  CPU_W_HDL_R_0_USER_RA_TRP1_6;
input  CPU_W_HDL_R_0_USER_RA_TRP1_7;
input  CPU_W_HDL_R_0_USER_RA_TRP1_9;
input  CPU_W_HDL_R_0_USER_REN_TRP1;
input  OSC_0_XTLOSC_O2F;
input  Glue_Logic_0_USER_WEN_TRP1;

    wire VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    RAM1K18 test_4463andcpuopration_COREEDAC_0_actram_R0C0 (.A_DOUT({
        nc0, nc1, nc2, nc3, nc4, CODE_FROM_RAM[12], CODE_FROM_RAM[11], 
        CODE_FROM_RAM[10], CODE_FROM_RAM[9], CODE_FROM_RAM[8], 
        CODE_FROM_RAM[7], CODE_FROM_RAM[6], CODE_FROM_RAM[5], 
        CODE_FROM_RAM[4], CODE_FROM_RAM[3], CODE_FROM_RAM[2], 
        CODE_FROM_RAM[1], CODE_FROM_RAM[0]}), .B_DOUT({nc5, nc6, nc7, 
        nc8, nc9, nc10, nc11, nc12, nc13, nc14, nc15, nc16, nc17, nc18, 
        nc19, nc20, nc21, nc22}), .BUSY(), .A_CLK(
        Bit_Count_16dec_i_1[3]), .A_DOUT_CLK(VCC_net_1), .A_ARST_N(
        VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({
        CPU_W_HDL_R_0_USER_REN_TRP1, VCC_net_1, VCC_net_1}), 
        .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({
        CPU_W_HDL_R_0_USER_RA_TRP1_9, GND_net_1, 
        CPU_W_HDL_R_0_USER_RA_TRP1_7, CPU_W_HDL_R_0_USER_RA_TRP1_6, 
        CPU_W_HDL_R_0_USER_RA_TRP1_5, CPU_W_HDL_R_0_USER_RA_TRP1_4, 
        CPU_W_HDL_R_0_USER_RA_TRP1_3, CPU_W_HDL_R_0_USER_RA_TRP1_2, 
        CPU_W_HDL_R_0_USER_RA_TRP1_1, CPU_W_HDL_R_0_USER_RA_TRP1_0, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .A_WEN({
        GND_net_1, GND_net_1}), .B_CLK(OSC_0_XTLOSC_O2F), .B_DOUT_CLK(
        VCC_net_1), .B_ARST_N(VCC_net_1), .B_DOUT_EN(VCC_net_1), 
        .B_BLK({Glue_Logic_0_USER_WEN_TRP1, VCC_net_1, VCC_net_1}), 
        .B_DOUT_ARST_N(GND_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        Glue_Logic_0_MSG_TRP1[7], Glue_Logic_0_MSG_TRP1[6], 
        Glue_Logic_0_MSG_TRP1[5], Glue_Logic_0_MSG_TRP1[4], 
        Glue_Logic_0_MSG_TRP1[3], Glue_Logic_0_MSG_TRP1[2], 
        Glue_Logic_0_MSG_TRP1[1], Glue_Logic_0_MSG_TRP1[0], CODED[4], 
        CODED[3], CODED[2], CODED[1], CODED[0]}), .B_ADDR({
        Glue_Logic_0_MSG_WA_TRP1[9], Glue_Logic_0_MSG_WA_TRP1[8], 
        Glue_Logic_0_MSG_WA_TRP1[7], Glue_Logic_0_MSG_WA_TRP1[6], 
        Glue_Logic_0_MSG_WA_TRP1[5], Glue_Logic_0_MSG_WA_TRP1[4], 
        Glue_Logic_0_MSG_WA_TRP1[3], Glue_Logic_0_MSG_WA_TRP1[2], 
        Glue_Logic_0_MSG_WA_TRP1[1], Glue_Logic_0_MSG_WA_TRP1[0], 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .B_WEN({
        VCC_net_1, VCC_net_1}), .A_EN(VCC_net_1), .A_DOUT_LAT(
        VCC_net_1), .A_WIDTH({VCC_net_1, GND_net_1, GND_net_1}), 
        .A_WMODE(GND_net_1), .B_EN(VCC_net_1), .B_DOUT_LAT(VCC_net_1), 
        .B_WIDTH({VCC_net_1, GND_net_1, GND_net_1}), .B_WMODE(
        GND_net_1), .SII_LOCK(GND_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_5(
       synd_w,
       CODE_FROM_RAM_9,
       CODE_FROM_RAM_7,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_6,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_4
    );
output [1:1] synd_w;
input  CODE_FROM_RAM_9;
input  CODE_FROM_RAM_7;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_6;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_4;

    wire \outp_3[0]_net_1 , GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_3[0]  (.A(CODE_FROM_RAM_9), .B(
        CODE_FROM_RAM_7), .C(CODE_FROM_RAM_11), .D(CODE_FROM_RAM_6), 
        .Y(\outp_3[0]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h96) )  \outp[0]  (.A(CODE_FROM_RAM_0), .B(
        CODE_FROM_RAM_4), .C(\outp_3[0]_net_1 ), .Y(synd_w[1]));
    
endmodule


module wide_xor_6s_3s_4294967295_4294967295_2s_4_0(
       synd_w,
       CODE_FROM_RAM_9,
       CODE_FROM_RAM_7,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_6,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_4
    );
output [1:1] synd_w;
input  CODE_FROM_RAM_9;
input  CODE_FROM_RAM_7;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_6;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_4;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    layer_xor_1s_3s_0_3s_1s_5 \genXOR[1].layer_xor_0  (.synd_w({
        synd_w[1]}), .CODE_FROM_RAM_9(CODE_FROM_RAM_9), 
        .CODE_FROM_RAM_7(CODE_FROM_RAM_7), .CODE_FROM_RAM_11(
        CODE_FROM_RAM_11), .CODE_FROM_RAM_6(CODE_FROM_RAM_6), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM_0), .CODE_FROM_RAM_4(
        CODE_FROM_RAM_4));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_8(
       outp_1_0,
       CODE_FROM_RAM_2,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_7,
       CODE_FROM_RAM_8,
       CODE_FROM_RAM_3,
       CODE_FROM_RAM_5,
       CODE_FROM_RAM_4,
       synd_w_4,
       synd_w_1,
       synd_w_2,
       synd_w_0,
       CPU_W_HDL_R_0_DataO_5,
       CPU_W_HDL_R_0_DataO_4,
       CPU_W_HDL_R_0_DataO_2,
       CPU_W_HDL_R_0_DataO_0,
       N_18,
       N_16,
       N_44,
       N_34_mux,
       m9_out,
       m4_out
    );
input  [0:0] outp_1_0;
input  CODE_FROM_RAM_2;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_7;
input  CODE_FROM_RAM_8;
input  CODE_FROM_RAM_3;
input  CODE_FROM_RAM_5;
input  CODE_FROM_RAM_4;
output synd_w_4;
input  synd_w_1;
input  synd_w_2;
input  synd_w_0;
output CPU_W_HDL_R_0_DataO_5;
output CPU_W_HDL_R_0_DataO_4;
output CPU_W_HDL_R_0_DataO_2;
output CPU_W_HDL_R_0_DataO_0;
output N_18;
output N_16;
output N_44;
output N_34_mux;
output m9_out;
output m4_out;

    wire \outp_1[0]_net_1 , GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h0090) )  \outp_RNIDUE71_1[0]  (.A(N_16), .B(
        outp_1_0[0]), .C(synd_w_4), .D(synd_w_1), .Y(m4_out));
    CFG4 #( .INIT(16'h9AAA) )  \outp_RNIO3J12_2[0]  (.A(
        CODE_FROM_RAM_8), .B(synd_w_0), .C(synd_w_2), .D(N_44), .Y(
        CPU_W_HDL_R_0_DataO_5));
    CFG4 #( .INIT(16'h9669) )  \outp[0]  (.A(CODE_FROM_RAM_4), .B(
        CODE_FROM_RAM_5), .C(N_18), .D(\outp_1[0]_net_1 ), .Y(synd_w_4)
        );
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h9) )  m17 (.A(CODE_FROM_RAM_7), .B(
        CODE_FROM_RAM_8), .Y(N_18));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h9) )  m15 (.A(CODE_FROM_RAM_3), .B(
        CODE_FROM_RAM_5), .Y(N_16));
    CFG4 #( .INIT(16'h6000) )  m11 (.A(outp_1_0[0]), .B(N_16), .C(
        synd_w_2), .D(synd_w_0), .Y(N_34_mux));
    CFG4 #( .INIT(16'hA6AA) )  \outp_RNIO3J12[0]  (.A(CODE_FROM_RAM_7), 
        .B(synd_w_4), .C(synd_w_1), .D(N_34_mux), .Y(
        CPU_W_HDL_R_0_DataO_4));
    CFG2 #( .INIT(4'h6) )  \outp_1[0]  (.A(CODE_FROM_RAM_2), .B(
        CODE_FROM_RAM_0), .Y(\outp_1[0]_net_1 ));
    CFG4 #( .INIT(16'h9AAA) )  \outp_RNIO3J12_0[0]  (.A(
        CODE_FROM_RAM_5), .B(synd_w_0), .C(synd_w_2), .D(m4_out), .Y(
        CPU_W_HDL_R_0_DataO_2));
    CFG4 #( .INIT(16'h6000) )  \outp_RNIDUE71[0]  (.A(N_16), .B(
        outp_1_0[0]), .C(synd_w_4), .D(synd_w_1), .Y(N_44));
    CFG4 #( .INIT(16'h9AAA) )  \outp_RNIO3J12_1[0]  (.A(
        CODE_FROM_RAM_3), .B(synd_w_0), .C(synd_w_2), .D(m9_out), .Y(
        CPU_W_HDL_R_0_DataO_0));
    CFG4 #( .INIT(16'h0900) )  \outp_RNIDUE71_0[0]  (.A(N_16), .B(
        outp_1_0[0]), .C(synd_w_4), .D(synd_w_1), .Y(m9_out));
    
endmodule


module wide_xor_6s_3s_4294967295_4294967295_2s_4_3(
       outp_1,
       CODE_FROM_RAM_2,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_7,
       CODE_FROM_RAM_8,
       CODE_FROM_RAM_3,
       CODE_FROM_RAM_5,
       CODE_FROM_RAM_4,
       synd_w_4,
       synd_w_1,
       synd_w_2,
       synd_w_0,
       CPU_W_HDL_R_0_DataO_5,
       CPU_W_HDL_R_0_DataO_4,
       CPU_W_HDL_R_0_DataO_2,
       CPU_W_HDL_R_0_DataO_0,
       N_18,
       N_16,
       N_44,
       N_34_mux,
       m9_out,
       m4_out
    );
input  [0:0] outp_1;
input  CODE_FROM_RAM_2;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_7;
input  CODE_FROM_RAM_8;
input  CODE_FROM_RAM_3;
input  CODE_FROM_RAM_5;
input  CODE_FROM_RAM_4;
output synd_w_4;
input  synd_w_1;
input  synd_w_2;
input  synd_w_0;
output CPU_W_HDL_R_0_DataO_5;
output CPU_W_HDL_R_0_DataO_4;
output CPU_W_HDL_R_0_DataO_2;
output CPU_W_HDL_R_0_DataO_0;
output N_18;
output N_16;
output N_44;
output N_34_mux;
output m9_out;
output m4_out;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    layer_xor_1s_3s_0_3s_1s_8 \genXOR[1].layer_xor_0  (.outp_1_0({
        outp_1[0]}), .CODE_FROM_RAM_2(CODE_FROM_RAM_2), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM_0), .CODE_FROM_RAM_7(
        CODE_FROM_RAM_7), .CODE_FROM_RAM_8(CODE_FROM_RAM_8), 
        .CODE_FROM_RAM_3(CODE_FROM_RAM_3), .CODE_FROM_RAM_5(
        CODE_FROM_RAM_5), .CODE_FROM_RAM_4(CODE_FROM_RAM_4), .synd_w_4(
        synd_w_4), .synd_w_1(synd_w_1), .synd_w_2(synd_w_2), .synd_w_0(
        synd_w_0), .CPU_W_HDL_R_0_DataO_5(CPU_W_HDL_R_0_DataO_5), 
        .CPU_W_HDL_R_0_DataO_4(CPU_W_HDL_R_0_DataO_4), 
        .CPU_W_HDL_R_0_DataO_2(CPU_W_HDL_R_0_DataO_2), 
        .CPU_W_HDL_R_0_DataO_0(CPU_W_HDL_R_0_DataO_0), .N_18(N_18), 
        .N_16(N_16), .N_44(N_44), .N_34_mux(N_34_mux), .m9_out(m9_out), 
        .m4_out(m4_out));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_7(
       outp_1,
       CODE_FROM_RAM_3,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_7
    );
output [0:0] outp_1;
input  CODE_FROM_RAM_3;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_7;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h96) )  \outp_1[0]  (.A(CODE_FROM_RAM_3), .B(
        CODE_FROM_RAM_0), .C(CODE_FROM_RAM_7), .Y(outp_1[0]));
    
endmodule


module wide_xor_6s_3s_4294967295_4294967295_2s_4_2(
       outp_1,
       CODE_FROM_RAM_3,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_7
    );
output [0:0] outp_1;
input  CODE_FROM_RAM_3;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_7;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    layer_xor_1s_3s_0_3s_1s_7 \genXOR[1].layer_xor_0  (.outp_1({
        outp_1[0]}), .CODE_FROM_RAM_3(CODE_FROM_RAM_3), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM_0), .CODE_FROM_RAM_7(
        CODE_FROM_RAM_7));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_4(
       synd_w,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_10,
       CODE_FROM_RAM_8,
       CODE_FROM_RAM_6,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_5
    );
output [0:0] synd_w;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_10;
input  CODE_FROM_RAM_8;
input  CODE_FROM_RAM_6;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_5;

    wire \outp_3[0]_net_1 , GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp_3[0]  (.A(CODE_FROM_RAM_11), .B(
        CODE_FROM_RAM_10), .C(CODE_FROM_RAM_8), .D(CODE_FROM_RAM_6), 
        .Y(\outp_3[0]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h96) )  \outp[0]  (.A(CODE_FROM_RAM_0), .B(
        CODE_FROM_RAM_5), .C(\outp_3[0]_net_1 ), .Y(synd_w[0]));
    
endmodule


module wide_xor_6s_3s_4294967295_4294967295_2s_4(
       synd_w,
       CODE_FROM_RAM_11,
       CODE_FROM_RAM_10,
       CODE_FROM_RAM_8,
       CODE_FROM_RAM_6,
       CODE_FROM_RAM_0,
       CODE_FROM_RAM_5
    );
output [0:0] synd_w;
input  CODE_FROM_RAM_11;
input  CODE_FROM_RAM_10;
input  CODE_FROM_RAM_8;
input  CODE_FROM_RAM_6;
input  CODE_FROM_RAM_0;
input  CODE_FROM_RAM_5;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    layer_xor_1s_3s_0_3s_1s_4 \genXOR[1].layer_xor_0  (.synd_w({
        synd_w[0]}), .CODE_FROM_RAM_11(CODE_FROM_RAM_11), 
        .CODE_FROM_RAM_10(CODE_FROM_RAM_10), .CODE_FROM_RAM_8(
        CODE_FROM_RAM_8), .CODE_FROM_RAM_6(CODE_FROM_RAM_6), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM_0), .CODE_FROM_RAM_5(
        CODE_FROM_RAM_5));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_6(
       synd_w,
       CODE_FROM_RAM_3,
       CODE_FROM_RAM_0,
       N_16,
       N_18
    );
output [2:2] synd_w;
input  CODE_FROM_RAM_3;
input  CODE_FROM_RAM_0;
input  N_16;
input  N_18;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(CODE_FROM_RAM_3), .B(
        CODE_FROM_RAM_0), .C(N_16), .D(N_18), .Y(synd_w[2]));
    
endmodule


module wide_xor_6s_3s_4294967295_4294967295_2s_4_1(
       synd_w,
       CODE_FROM_RAM_3,
       CODE_FROM_RAM_0,
       N_16,
       N_18
    );
output [2:2] synd_w;
input  CODE_FROM_RAM_3;
input  CODE_FROM_RAM_0;
input  N_16;
input  N_18;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    layer_xor_1s_3s_0_3s_1s_6 \genXOR[1].layer_xor_0  (.synd_w({
        synd_w[2]}), .CODE_FROM_RAM_3(CODE_FROM_RAM_3), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM_0), .N_16(N_16), .N_18(N_18));
    
endmodule


module 
        test_4463andcpuopration_COREEDAC_0_ham_dec_vlog_8s_5_0_4294967295_4294967295_0(
        
       CODE_FROM_RAM,
       CPU_W_HDL_R_0_DataO
    );
input  [12:0] CODE_FROM_RAM;
output [7:0] CPU_W_HDL_R_0_DataO;

    wire \synd_w[4] , \synd_w[1] , N_34_mux, \synd_w[0] , \synd_w[2] , 
        m4_out, N_44, m9_out, N_16, N_18, \outp_1[0] , GND_net_1, 
        VCC_net_1;
    
    CFG4 #( .INIT(16'hA6AA) )  \re_code[8]  (.A(CODE_FROM_RAM[8]), .B(
        \synd_w[0] ), .C(\synd_w[2] ), .D(N_44), .Y(
        CPU_W_HDL_R_0_DataO[3]));
    CFG4 #( .INIT(16'hA6AA) )  \re_code[6]  (.A(CODE_FROM_RAM[6]), .B(
        \synd_w[0] ), .C(\synd_w[2] ), .D(m4_out), .Y(
        CPU_W_HDL_R_0_DataO[1]));
    wide_xor_6s_3s_4294967295_4294967295_2s_4_0 wide_xor_1 (.synd_w({
        \synd_w[1] }), .CODE_FROM_RAM_9(CODE_FROM_RAM[10]), 
        .CODE_FROM_RAM_7(CODE_FROM_RAM[8]), .CODE_FROM_RAM_11(
        CODE_FROM_RAM[12]), .CODE_FROM_RAM_6(CODE_FROM_RAM[7]), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM[1]), .CODE_FROM_RAM_4(
        CODE_FROM_RAM[5]));
    GND GND (.Y(GND_net_1));
    wide_xor_6s_3s_4294967295_4294967295_2s_4_3 wide_xor_4 (.outp_1({
        \outp_1[0] }), .CODE_FROM_RAM_2(CODE_FROM_RAM[6]), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM[4]), .CODE_FROM_RAM_7(
        CODE_FROM_RAM[11]), .CODE_FROM_RAM_8(CODE_FROM_RAM[12]), 
        .CODE_FROM_RAM_3(CODE_FROM_RAM[7]), .CODE_FROM_RAM_5(
        CODE_FROM_RAM[9]), .CODE_FROM_RAM_4(CODE_FROM_RAM[8]), 
        .synd_w_4(\synd_w[4] ), .synd_w_1(\synd_w[1] ), .synd_w_2(
        \synd_w[2] ), .synd_w_0(\synd_w[0] ), .CPU_W_HDL_R_0_DataO_5(
        CPU_W_HDL_R_0_DataO[7]), .CPU_W_HDL_R_0_DataO_4(
        CPU_W_HDL_R_0_DataO[6]), .CPU_W_HDL_R_0_DataO_2(
        CPU_W_HDL_R_0_DataO[4]), .CPU_W_HDL_R_0_DataO_0(
        CPU_W_HDL_R_0_DataO[2]), .N_18(N_18), .N_16(N_16), .N_44(N_44), 
        .N_34_mux(N_34_mux), .m9_out(m9_out), .m4_out(m4_out));
    CFG4 #( .INIT(16'hA6AA) )  \re_code[10]  (.A(CODE_FROM_RAM[10]), 
        .B(\synd_w[0] ), .C(\synd_w[2] ), .D(m9_out), .Y(
        CPU_W_HDL_R_0_DataO[5]));
    VCC VCC (.Y(VCC_net_1));
    wide_xor_6s_3s_4294967295_4294967295_2s_4_2 wide_xor_3 (.outp_1({
        \outp_1[0] }), .CODE_FROM_RAM_3(CODE_FROM_RAM[6]), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM[3]), .CODE_FROM_RAM_7(
        CODE_FROM_RAM[10]));
    wide_xor_6s_3s_4294967295_4294967295_2s_4 wide_xor_0 (.synd_w({
        \synd_w[0] }), .CODE_FROM_RAM_11(CODE_FROM_RAM[11]), 
        .CODE_FROM_RAM_10(CODE_FROM_RAM[10]), .CODE_FROM_RAM_8(
        CODE_FROM_RAM[8]), .CODE_FROM_RAM_6(CODE_FROM_RAM[6]), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM[0]), .CODE_FROM_RAM_5(
        CODE_FROM_RAM[5]));
    CFG4 #( .INIT(16'h9AAA) )  \re_code[5]  (.A(CODE_FROM_RAM[5]), .B(
        \synd_w[4] ), .C(\synd_w[1] ), .D(N_34_mux), .Y(
        CPU_W_HDL_R_0_DataO[0]));
    wide_xor_6s_3s_4294967295_4294967295_2s_4_1 wide_xor_2 (.synd_w({
        \synd_w[2] }), .CODE_FROM_RAM_3(CODE_FROM_RAM[5]), 
        .CODE_FROM_RAM_0(CODE_FROM_RAM[2]), .N_16(N_16), .N_18(N_18));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_1(
       CODED_2,
       CODED,
       Glue_Logic_0_MSG_TRP1_7,
       Glue_Logic_0_MSG_TRP1_2,
       Glue_Logic_0_MSG_TRP1_0
    );
input  [4:4] CODED_2;
output [2:2] CODED;
input  Glue_Logic_0_MSG_TRP1_7;
input  Glue_Logic_0_MSG_TRP1_2;
input  Glue_Logic_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(Glue_Logic_0_MSG_TRP1_7), 
        .B(Glue_Logic_0_MSG_TRP1_2), .C(Glue_Logic_0_MSG_TRP1_0), .D(
        CODED_2[4]), .Y(CODED[2]));
    
endmodule


module wide_xor_5s_3s_4294967295_4294967295_2s_4_1(
       CODED_2,
       CODED,
       Glue_Logic_0_MSG_TRP1_7,
       Glue_Logic_0_MSG_TRP1_2,
       Glue_Logic_0_MSG_TRP1_0
    );
input  [4:4] CODED_2;
output [2:2] CODED;
input  Glue_Logic_0_MSG_TRP1_7;
input  Glue_Logic_0_MSG_TRP1_2;
input  Glue_Logic_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    layer_xor_1s_3s_0_3s_1s_1 \genXOR[1].layer_xor_0  (.CODED_2({
        CODED_2[4]}), .CODED({CODED[2]}), .Glue_Logic_0_MSG_TRP1_7(
        Glue_Logic_0_MSG_TRP1_7), .Glue_Logic_0_MSG_TRP1_2(
        Glue_Logic_0_MSG_TRP1_2), .Glue_Logic_0_MSG_TRP1_0(
        Glue_Logic_0_MSG_TRP1_0));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_0(
       CODED_2,
       CODED,
       Glue_Logic_0_MSG_TRP1_7,
       Glue_Logic_0_MSG_TRP1_2,
       Glue_Logic_0_MSG_TRP1_0
    );
input  [1:1] CODED_2;
output [1:1] CODED;
input  Glue_Logic_0_MSG_TRP1_7;
input  Glue_Logic_0_MSG_TRP1_2;
input  Glue_Logic_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(Glue_Logic_0_MSG_TRP1_7), 
        .B(Glue_Logic_0_MSG_TRP1_2), .C(Glue_Logic_0_MSG_TRP1_0), .D(
        CODED_2[1]), .Y(CODED[1]));
    
endmodule


module wide_xor_5s_3s_4294967295_4294967295_2s_4_0(
       CODED_2,
       CODED,
       Glue_Logic_0_MSG_TRP1_7,
       Glue_Logic_0_MSG_TRP1_2,
       Glue_Logic_0_MSG_TRP1_0
    );
input  [1:1] CODED_2;
output [1:1] CODED;
input  Glue_Logic_0_MSG_TRP1_7;
input  Glue_Logic_0_MSG_TRP1_2;
input  Glue_Logic_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    layer_xor_1s_3s_0_3s_1s_0 \genXOR[1].layer_xor_0  (.CODED_2({
        CODED_2[1]}), .CODED({CODED[1]}), .Glue_Logic_0_MSG_TRP1_7(
        Glue_Logic_0_MSG_TRP1_7), .Glue_Logic_0_MSG_TRP1_2(
        Glue_Logic_0_MSG_TRP1_2), .Glue_Logic_0_MSG_TRP1_0(
        Glue_Logic_0_MSG_TRP1_0));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_3(
       CODED_2,
       CODED,
       Glue_Logic_0_MSG_TRP1_3,
       Glue_Logic_0_MSG_TRP1_5,
       Glue_Logic_0_MSG_TRP1_6,
       Glue_Logic_0_MSG_TRP1_2,
       Glue_Logic_0_MSG_TRP1_0
    );
output [4:4] CODED_2;
output [4:4] CODED;
input  Glue_Logic_0_MSG_TRP1_3;
input  Glue_Logic_0_MSG_TRP1_5;
input  Glue_Logic_0_MSG_TRP1_6;
input  Glue_Logic_0_MSG_TRP1_2;
input  Glue_Logic_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h6) )  \outp_2[0]  (.A(Glue_Logic_0_MSG_TRP1_3), 
        .B(Glue_Logic_0_MSG_TRP1_5), .Y(CODED_2[4]));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(Glue_Logic_0_MSG_TRP1_6), 
        .B(Glue_Logic_0_MSG_TRP1_2), .C(CODED_2[4]), .D(
        Glue_Logic_0_MSG_TRP1_0), .Y(CODED[4]));
    
endmodule


module wide_xor_5s_3s_4294967295_4294967295_2s_4_3(
       CODED_2,
       CODED,
       Glue_Logic_0_MSG_TRP1_3,
       Glue_Logic_0_MSG_TRP1_5,
       Glue_Logic_0_MSG_TRP1_6,
       Glue_Logic_0_MSG_TRP1_2,
       Glue_Logic_0_MSG_TRP1_0
    );
output [4:4] CODED_2;
output [4:4] CODED;
input  Glue_Logic_0_MSG_TRP1_3;
input  Glue_Logic_0_MSG_TRP1_5;
input  Glue_Logic_0_MSG_TRP1_6;
input  Glue_Logic_0_MSG_TRP1_2;
input  Glue_Logic_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    layer_xor_1s_3s_0_3s_1s_3 \genXOR[1].layer_xor_0  (.CODED_2({
        CODED_2[4]}), .CODED({CODED[4]}), .Glue_Logic_0_MSG_TRP1_3(
        Glue_Logic_0_MSG_TRP1_3), .Glue_Logic_0_MSG_TRP1_5(
        Glue_Logic_0_MSG_TRP1_5), .Glue_Logic_0_MSG_TRP1_6(
        Glue_Logic_0_MSG_TRP1_6), .Glue_Logic_0_MSG_TRP1_2(
        Glue_Logic_0_MSG_TRP1_2), .Glue_Logic_0_MSG_TRP1_0(
        Glue_Logic_0_MSG_TRP1_0));
    
endmodule


module layer_xor_1s_3s_0_3s_1s(
       CODED_2,
       CODED,
       Glue_Logic_0_MSG_TRP1_3,
       Glue_Logic_0_MSG_TRP1_5,
       Glue_Logic_0_MSG_TRP1_6,
       Glue_Logic_0_MSG_TRP1_1,
       Glue_Logic_0_MSG_TRP1_0
    );
output [1:1] CODED_2;
output [0:0] CODED;
input  Glue_Logic_0_MSG_TRP1_3;
input  Glue_Logic_0_MSG_TRP1_5;
input  Glue_Logic_0_MSG_TRP1_6;
input  Glue_Logic_0_MSG_TRP1_1;
input  Glue_Logic_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG2 #( .INIT(4'h6) )  \outp_2[0]  (.A(Glue_Logic_0_MSG_TRP1_3), 
        .B(Glue_Logic_0_MSG_TRP1_5), .Y(CODED_2[1]));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(Glue_Logic_0_MSG_TRP1_6), 
        .B(Glue_Logic_0_MSG_TRP1_1), .C(Glue_Logic_0_MSG_TRP1_0), .D(
        CODED_2[1]), .Y(CODED[0]));
    
endmodule


module wide_xor_5s_3s_4294967295_4294967295_2s_4(
       CODED_2,
       CODED,
       Glue_Logic_0_MSG_TRP1_3,
       Glue_Logic_0_MSG_TRP1_5,
       Glue_Logic_0_MSG_TRP1_6,
       Glue_Logic_0_MSG_TRP1_1,
       Glue_Logic_0_MSG_TRP1_0
    );
output [1:1] CODED_2;
output [0:0] CODED;
input  Glue_Logic_0_MSG_TRP1_3;
input  Glue_Logic_0_MSG_TRP1_5;
input  Glue_Logic_0_MSG_TRP1_6;
input  Glue_Logic_0_MSG_TRP1_1;
input  Glue_Logic_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    layer_xor_1s_3s_0_3s_1s \genXOR[1].layer_xor_0  (.CODED_2({
        CODED_2[1]}), .CODED({CODED[0]}), .Glue_Logic_0_MSG_TRP1_3(
        Glue_Logic_0_MSG_TRP1_3), .Glue_Logic_0_MSG_TRP1_5(
        Glue_Logic_0_MSG_TRP1_5), .Glue_Logic_0_MSG_TRP1_6(
        Glue_Logic_0_MSG_TRP1_6), .Glue_Logic_0_MSG_TRP1_1(
        Glue_Logic_0_MSG_TRP1_1), .Glue_Logic_0_MSG_TRP1_0(
        Glue_Logic_0_MSG_TRP1_0));
    
endmodule


module layer_xor_1s_3s_0_3s_1s_2(
       CODED,
       Glue_Logic_0_MSG_TRP1_4,
       Glue_Logic_0_MSG_TRP1_3,
       Glue_Logic_0_MSG_TRP1_1,
       Glue_Logic_0_MSG_TRP1_0
    );
output [3:3] CODED;
input  Glue_Logic_0_MSG_TRP1_4;
input  Glue_Logic_0_MSG_TRP1_3;
input  Glue_Logic_0_MSG_TRP1_1;
input  Glue_Logic_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h6996) )  \outp[0]  (.A(Glue_Logic_0_MSG_TRP1_4), 
        .B(Glue_Logic_0_MSG_TRP1_3), .C(Glue_Logic_0_MSG_TRP1_1), .D(
        Glue_Logic_0_MSG_TRP1_0), .Y(CODED[3]));
    
endmodule


module wide_xor_5s_3s_4294967295_4294967295_2s_4_2(
       CODED,
       Glue_Logic_0_MSG_TRP1_4,
       Glue_Logic_0_MSG_TRP1_3,
       Glue_Logic_0_MSG_TRP1_1,
       Glue_Logic_0_MSG_TRP1_0
    );
output [3:3] CODED;
input  Glue_Logic_0_MSG_TRP1_4;
input  Glue_Logic_0_MSG_TRP1_3;
input  Glue_Logic_0_MSG_TRP1_1;
input  Glue_Logic_0_MSG_TRP1_0;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    layer_xor_1s_3s_0_3s_1s_2 \genXOR[1].layer_xor_0  (.CODED({
        CODED[3]}), .Glue_Logic_0_MSG_TRP1_4(Glue_Logic_0_MSG_TRP1_4), 
        .Glue_Logic_0_MSG_TRP1_3(Glue_Logic_0_MSG_TRP1_3), 
        .Glue_Logic_0_MSG_TRP1_1(Glue_Logic_0_MSG_TRP1_1), 
        .Glue_Logic_0_MSG_TRP1_0(Glue_Logic_0_MSG_TRP1_0));
    
endmodule


module 
        test_4463andcpuopration_COREEDAC_0_ham_enc_vlog_8s_5_4294967295_4294967295(
        
       Glue_Logic_0_MSG_TRP1,
       CODED
    );
input  [7:0] Glue_Logic_0_MSG_TRP1;
output [4:0] CODED;

    wire \CODED_2[1] , \CODED_2[4] , GND_net_1, VCC_net_1;
    
    wide_xor_5s_3s_4294967295_4294967295_2s_4_1 wide_xor_2 (.CODED_2({
        \CODED_2[4] }), .CODED({CODED[2]}), .Glue_Logic_0_MSG_TRP1_7(
        Glue_Logic_0_MSG_TRP1[7]), .Glue_Logic_0_MSG_TRP1_2(
        Glue_Logic_0_MSG_TRP1[2]), .Glue_Logic_0_MSG_TRP1_0(
        Glue_Logic_0_MSG_TRP1[0]));
    wide_xor_5s_3s_4294967295_4294967295_2s_4_0 wide_xor_1 (.CODED_2({
        \CODED_2[1] }), .CODED({CODED[1]}), .Glue_Logic_0_MSG_TRP1_7(
        Glue_Logic_0_MSG_TRP1[7]), .Glue_Logic_0_MSG_TRP1_2(
        Glue_Logic_0_MSG_TRP1[2]), .Glue_Logic_0_MSG_TRP1_0(
        Glue_Logic_0_MSG_TRP1[0]));
    wide_xor_5s_3s_4294967295_4294967295_2s_4_3 wide_xor_4 (.CODED_2({
        \CODED_2[4] }), .CODED({CODED[4]}), .Glue_Logic_0_MSG_TRP1_3(
        Glue_Logic_0_MSG_TRP1[4]), .Glue_Logic_0_MSG_TRP1_5(
        Glue_Logic_0_MSG_TRP1[6]), .Glue_Logic_0_MSG_TRP1_6(
        Glue_Logic_0_MSG_TRP1[7]), .Glue_Logic_0_MSG_TRP1_2(
        Glue_Logic_0_MSG_TRP1[3]), .Glue_Logic_0_MSG_TRP1_0(
        Glue_Logic_0_MSG_TRP1[1]));
    VCC VCC (.Y(VCC_net_1));
    wide_xor_5s_3s_4294967295_4294967295_2s_4 wide_xor_0 (.CODED_2({
        \CODED_2[1] }), .CODED({CODED[0]}), .Glue_Logic_0_MSG_TRP1_3(
        Glue_Logic_0_MSG_TRP1[3]), .Glue_Logic_0_MSG_TRP1_5(
        Glue_Logic_0_MSG_TRP1[5]), .Glue_Logic_0_MSG_TRP1_6(
        Glue_Logic_0_MSG_TRP1[6]), .Glue_Logic_0_MSG_TRP1_1(
        Glue_Logic_0_MSG_TRP1[1]), .Glue_Logic_0_MSG_TRP1_0(
        Glue_Logic_0_MSG_TRP1[0]));
    GND GND (.Y(GND_net_1));
    wide_xor_5s_3s_4294967295_4294967295_2s_4_2 wide_xor_3 (.CODED({
        CODED[3]}), .Glue_Logic_0_MSG_TRP1_4(Glue_Logic_0_MSG_TRP1[5]), 
        .Glue_Logic_0_MSG_TRP1_3(Glue_Logic_0_MSG_TRP1[4]), 
        .Glue_Logic_0_MSG_TRP1_1(Glue_Logic_0_MSG_TRP1[2]), 
        .Glue_Logic_0_MSG_TRP1_0(Glue_Logic_0_MSG_TRP1[1]));
    
endmodule


module test_4463andcpuopration_COREEDAC_0_ecc_Z2(
       Glue_Logic_0_MSG_TRP1,
       CODED,
       CODE_FROM_RAM,
       CPU_W_HDL_R_0_DataO
    );
input  [7:0] Glue_Logic_0_MSG_TRP1;
output [4:0] CODED;
input  [12:0] CODE_FROM_RAM;
output [7:0] CPU_W_HDL_R_0_DataO;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    
        test_4463andcpuopration_COREEDAC_0_ham_dec_vlog_8s_5_0_4294967295_4294967295_0 
        test_4463andcpuopration_COREEDAC_0_decoder_0 (.CODE_FROM_RAM({
        CODE_FROM_RAM[12], CODE_FROM_RAM[11], CODE_FROM_RAM[10], 
        CODE_FROM_RAM[9], CODE_FROM_RAM[8], CODE_FROM_RAM[7], 
        CODE_FROM_RAM[6], CODE_FROM_RAM[5], CODE_FROM_RAM[4], 
        CODE_FROM_RAM[3], CODE_FROM_RAM[2], CODE_FROM_RAM[1], 
        CODE_FROM_RAM[0]}), .CPU_W_HDL_R_0_DataO({
        CPU_W_HDL_R_0_DataO[7], CPU_W_HDL_R_0_DataO[6], 
        CPU_W_HDL_R_0_DataO[5], CPU_W_HDL_R_0_DataO[4], 
        CPU_W_HDL_R_0_DataO[3], CPU_W_HDL_R_0_DataO[2], 
        CPU_W_HDL_R_0_DataO[1], CPU_W_HDL_R_0_DataO[0]}));
    
        test_4463andcpuopration_COREEDAC_0_ham_enc_vlog_8s_5_4294967295_4294967295 
        test_4463andcpuopration_COREEDAC_0_encoder_0 (
        .Glue_Logic_0_MSG_TRP1({Glue_Logic_0_MSG_TRP1[7], 
        Glue_Logic_0_MSG_TRP1[6], Glue_Logic_0_MSG_TRP1[5], 
        Glue_Logic_0_MSG_TRP1[4], Glue_Logic_0_MSG_TRP1[3], 
        Glue_Logic_0_MSG_TRP1[2], Glue_Logic_0_MSG_TRP1[1], 
        Glue_Logic_0_MSG_TRP1[0]}), .CODED({CODED[4], CODED[3], 
        CODED[2], CODED[1], CODED[0]}));
    GND GND (.Y(GND_net_1));
    
endmodule


module test_4463andcpuopration_COREEDAC_0_sub_edac_Z3(
       Glue_Logic_0_MSG_TRP1,
       CODED,
       CODE_FROM_RAM,
       CPU_W_HDL_R_0_DataO
    );
input  [7:0] Glue_Logic_0_MSG_TRP1;
output [4:0] CODED;
input  [12:0] CODE_FROM_RAM;
output [7:0] CPU_W_HDL_R_0_DataO;

    wire GND_net_1, VCC_net_1;
    
    test_4463andcpuopration_COREEDAC_0_ecc_Z2 
        test_4463andcpuopration_COREEDAC_0_ecc_0 (
        .Glue_Logic_0_MSG_TRP1({Glue_Logic_0_MSG_TRP1[7], 
        Glue_Logic_0_MSG_TRP1[6], Glue_Logic_0_MSG_TRP1[5], 
        Glue_Logic_0_MSG_TRP1[4], Glue_Logic_0_MSG_TRP1[3], 
        Glue_Logic_0_MSG_TRP1[2], Glue_Logic_0_MSG_TRP1[1], 
        Glue_Logic_0_MSG_TRP1[0]}), .CODED({CODED[4], CODED[3], 
        CODED[2], CODED[1], CODED[0]}), .CODE_FROM_RAM({
        CODE_FROM_RAM[12], CODE_FROM_RAM[11], CODE_FROM_RAM[10], 
        CODE_FROM_RAM[9], CODE_FROM_RAM[8], CODE_FROM_RAM[7], 
        CODE_FROM_RAM[6], CODE_FROM_RAM[5], CODE_FROM_RAM[4], 
        CODE_FROM_RAM[3], CODE_FROM_RAM[2], CODE_FROM_RAM[1], 
        CODE_FROM_RAM[0]}), .CPU_W_HDL_R_0_DataO({
        CPU_W_HDL_R_0_DataO[7], CPU_W_HDL_R_0_DataO[6], 
        CPU_W_HDL_R_0_DataO[5], CPU_W_HDL_R_0_DataO[4], 
        CPU_W_HDL_R_0_DataO[3], CPU_W_HDL_R_0_DataO[2], 
        CPU_W_HDL_R_0_DataO[1], CPU_W_HDL_R_0_DataO[0]}));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module test_4463andcpuopration_COREEDAC_0_edac_Z4(
       Glue_Logic_0_MSG_TRP1,
       CODED,
       CODE_FROM_RAM,
       CPU_W_HDL_R_0_DataO
    );
input  [7:0] Glue_Logic_0_MSG_TRP1;
output [4:0] CODED;
input  [12:0] CODE_FROM_RAM;
output [7:0] CPU_W_HDL_R_0_DataO;

    wire GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    test_4463andcpuopration_COREEDAC_0_sub_edac_Z3 
        test_4463andcpuopration_COREEDAC_0_sub_edac_0 (
        .Glue_Logic_0_MSG_TRP1({Glue_Logic_0_MSG_TRP1[7], 
        Glue_Logic_0_MSG_TRP1[6], Glue_Logic_0_MSG_TRP1[5], 
        Glue_Logic_0_MSG_TRP1[4], Glue_Logic_0_MSG_TRP1[3], 
        Glue_Logic_0_MSG_TRP1[2], Glue_Logic_0_MSG_TRP1[1], 
        Glue_Logic_0_MSG_TRP1[0]}), .CODED({CODED[4], CODED[3], 
        CODED[2], CODED[1], CODED[0]}), .CODE_FROM_RAM({
        CODE_FROM_RAM[12], CODE_FROM_RAM[11], CODE_FROM_RAM[10], 
        CODE_FROM_RAM[9], CODE_FROM_RAM[8], CODE_FROM_RAM[7], 
        CODE_FROM_RAM[6], CODE_FROM_RAM[5], CODE_FROM_RAM[4], 
        CODE_FROM_RAM[3], CODE_FROM_RAM[2], CODE_FROM_RAM[1], 
        CODE_FROM_RAM[0]}), .CPU_W_HDL_R_0_DataO({
        CPU_W_HDL_R_0_DataO[7], CPU_W_HDL_R_0_DataO[6], 
        CPU_W_HDL_R_0_DataO[5], CPU_W_HDL_R_0_DataO[4], 
        CPU_W_HDL_R_0_DataO[3], CPU_W_HDL_R_0_DataO[2], 
        CPU_W_HDL_R_0_DataO[1], CPU_W_HDL_R_0_DataO[0]}));
    GND GND (.Y(GND_net_1));
    
endmodule


module test_4463andcpuopration_COREEDAC_0_COREEDAC_Z5(
       Glue_Logic_0_MSG_TRP1,
       CPU_W_HDL_R_0_DataO,
       Bit_Count_16dec_i_1,
       Glue_Logic_0_MSG_WA_TRP1,
       CPU_W_HDL_R_0_USER_RA_TRP1_0,
       CPU_W_HDL_R_0_USER_RA_TRP1_1,
       CPU_W_HDL_R_0_USER_RA_TRP1_2,
       CPU_W_HDL_R_0_USER_RA_TRP1_3,
       CPU_W_HDL_R_0_USER_RA_TRP1_4,
       CPU_W_HDL_R_0_USER_RA_TRP1_5,
       CPU_W_HDL_R_0_USER_RA_TRP1_6,
       CPU_W_HDL_R_0_USER_RA_TRP1_7,
       CPU_W_HDL_R_0_USER_RA_TRP1_9,
       CPU_W_HDL_R_0_USER_REN_TRP1,
       OSC_0_XTLOSC_O2F,
       Glue_Logic_0_USER_WEN_TRP1
    );
input  [7:0] Glue_Logic_0_MSG_TRP1;
output [7:0] CPU_W_HDL_R_0_DataO;
input  [3:3] Bit_Count_16dec_i_1;
input  [9:0] Glue_Logic_0_MSG_WA_TRP1;
input  CPU_W_HDL_R_0_USER_RA_TRP1_0;
input  CPU_W_HDL_R_0_USER_RA_TRP1_1;
input  CPU_W_HDL_R_0_USER_RA_TRP1_2;
input  CPU_W_HDL_R_0_USER_RA_TRP1_3;
input  CPU_W_HDL_R_0_USER_RA_TRP1_4;
input  CPU_W_HDL_R_0_USER_RA_TRP1_5;
input  CPU_W_HDL_R_0_USER_RA_TRP1_6;
input  CPU_W_HDL_R_0_USER_RA_TRP1_7;
input  CPU_W_HDL_R_0_USER_RA_TRP1_9;
input  CPU_W_HDL_R_0_USER_REN_TRP1;
input  OSC_0_XTLOSC_O2F;
input  Glue_Logic_0_USER_WEN_TRP1;

    wire \CODED[0] , \CODED[1] , \CODED[2] , \CODED[3] , \CODED[4] , 
        \CODE_FROM_RAM[0] , \CODE_FROM_RAM[1] , \CODE_FROM_RAM[2] , 
        \CODE_FROM_RAM[3] , \CODE_FROM_RAM[4] , \CODE_FROM_RAM[5] , 
        \CODE_FROM_RAM[6] , \CODE_FROM_RAM[7] , \CODE_FROM_RAM[8] , 
        \CODE_FROM_RAM[9] , \CODE_FROM_RAM[10] , \CODE_FROM_RAM[11] , 
        \CODE_FROM_RAM[12] , GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    test_4463andcpuopration_COREEDAC_0_actram 
        \lsram_g4.test_4463andcpuopration_COREEDAC_0_actram_0  (
        .CODE_FROM_RAM({\CODE_FROM_RAM[12] , \CODE_FROM_RAM[11] , 
        \CODE_FROM_RAM[10] , \CODE_FROM_RAM[9] , \CODE_FROM_RAM[8] , 
        \CODE_FROM_RAM[7] , \CODE_FROM_RAM[6] , \CODE_FROM_RAM[5] , 
        \CODE_FROM_RAM[4] , \CODE_FROM_RAM[3] , \CODE_FROM_RAM[2] , 
        \CODE_FROM_RAM[1] , \CODE_FROM_RAM[0] }), .Bit_Count_16dec_i_1({
        Bit_Count_16dec_i_1[3]}), .CODED({\CODED[4] , \CODED[3] , 
        \CODED[2] , \CODED[1] , \CODED[0] }), .Glue_Logic_0_MSG_TRP1({
        Glue_Logic_0_MSG_TRP1[7], Glue_Logic_0_MSG_TRP1[6], 
        Glue_Logic_0_MSG_TRP1[5], Glue_Logic_0_MSG_TRP1[4], 
        Glue_Logic_0_MSG_TRP1[3], Glue_Logic_0_MSG_TRP1[2], 
        Glue_Logic_0_MSG_TRP1[1], Glue_Logic_0_MSG_TRP1[0]}), 
        .Glue_Logic_0_MSG_WA_TRP1({Glue_Logic_0_MSG_WA_TRP1[9], 
        Glue_Logic_0_MSG_WA_TRP1[8], Glue_Logic_0_MSG_WA_TRP1[7], 
        Glue_Logic_0_MSG_WA_TRP1[6], Glue_Logic_0_MSG_WA_TRP1[5], 
        Glue_Logic_0_MSG_WA_TRP1[4], Glue_Logic_0_MSG_WA_TRP1[3], 
        Glue_Logic_0_MSG_WA_TRP1[2], Glue_Logic_0_MSG_WA_TRP1[1], 
        Glue_Logic_0_MSG_WA_TRP1[0]}), .CPU_W_HDL_R_0_USER_RA_TRP1_0(
        CPU_W_HDL_R_0_USER_RA_TRP1_0), .CPU_W_HDL_R_0_USER_RA_TRP1_1(
        CPU_W_HDL_R_0_USER_RA_TRP1_1), .CPU_W_HDL_R_0_USER_RA_TRP1_2(
        CPU_W_HDL_R_0_USER_RA_TRP1_2), .CPU_W_HDL_R_0_USER_RA_TRP1_3(
        CPU_W_HDL_R_0_USER_RA_TRP1_3), .CPU_W_HDL_R_0_USER_RA_TRP1_4(
        CPU_W_HDL_R_0_USER_RA_TRP1_4), .CPU_W_HDL_R_0_USER_RA_TRP1_5(
        CPU_W_HDL_R_0_USER_RA_TRP1_5), .CPU_W_HDL_R_0_USER_RA_TRP1_6(
        CPU_W_HDL_R_0_USER_RA_TRP1_6), .CPU_W_HDL_R_0_USER_RA_TRP1_7(
        CPU_W_HDL_R_0_USER_RA_TRP1_7), .CPU_W_HDL_R_0_USER_RA_TRP1_9(
        CPU_W_HDL_R_0_USER_RA_TRP1_9), .CPU_W_HDL_R_0_USER_REN_TRP1(
        CPU_W_HDL_R_0_USER_REN_TRP1), .OSC_0_XTLOSC_O2F(
        OSC_0_XTLOSC_O2F), .Glue_Logic_0_USER_WEN_TRP1(
        Glue_Logic_0_USER_WEN_TRP1));
    test_4463andcpuopration_COREEDAC_0_edac_Z4 
        test_4463andcpuopration_COREEDAC_0_edac_0 (
        .Glue_Logic_0_MSG_TRP1({Glue_Logic_0_MSG_TRP1[7], 
        Glue_Logic_0_MSG_TRP1[6], Glue_Logic_0_MSG_TRP1[5], 
        Glue_Logic_0_MSG_TRP1[4], Glue_Logic_0_MSG_TRP1[3], 
        Glue_Logic_0_MSG_TRP1[2], Glue_Logic_0_MSG_TRP1[1], 
        Glue_Logic_0_MSG_TRP1[0]}), .CODED({\CODED[4] , \CODED[3] , 
        \CODED[2] , \CODED[1] , \CODED[0] }), .CODE_FROM_RAM({
        \CODE_FROM_RAM[12] , \CODE_FROM_RAM[11] , \CODE_FROM_RAM[10] , 
        \CODE_FROM_RAM[9] , \CODE_FROM_RAM[8] , \CODE_FROM_RAM[7] , 
        \CODE_FROM_RAM[6] , \CODE_FROM_RAM[5] , \CODE_FROM_RAM[4] , 
        \CODE_FROM_RAM[3] , \CODE_FROM_RAM[2] , \CODE_FROM_RAM[1] , 
        \CODE_FROM_RAM[0] }), .CPU_W_HDL_R_0_DataO({
        CPU_W_HDL_R_0_DataO[7], CPU_W_HDL_R_0_DataO[6], 
        CPU_W_HDL_R_0_DataO[5], CPU_W_HDL_R_0_DataO[4], 
        CPU_W_HDL_R_0_DataO[3], CPU_W_HDL_R_0_DataO[2], 
        CPU_W_HDL_R_0_DataO[1], CPU_W_HDL_R_0_DataO[0]}));
    GND GND (.Y(GND_net_1));
    
endmodule


module RSControl(
       Bit_Count_16dec_i_1,
       RSControl_0_DATAINP,
       CPU_W_HDL_R_0_DataO,
       RSControl_0_NGRST,
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       RSControl_0_START,
       TM_RSENC_0_RFD,
       ENCRC,
       TM_RSENC_0_RFS
    );
input  [3:3] Bit_Count_16dec_i_1;
output [7:0] RSControl_0_DATAINP;
input  [7:0] CPU_W_HDL_R_0_DataO;
output RSControl_0_NGRST;
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
output RSControl_0_START;
input  TM_RSENC_0_RFD;
input  ENCRC;
input  TM_RSENC_0_RFS;

    wire NGRST_net_1, \Data_Buff[1]_net_1 , VCC_net_1, N_75_i_0, 
        GND_net_1, \Data_Buff[2]_net_1 , \Data_Buff[3]_net_1 , 
        \Data_Buff[4]_net_1 , \Data_Buff[5]_net_1 , 
        \Data_Buff[6]_net_1 , \Data_Buff[7]_net_1 , 
        \Data_Buff[0]_net_1 , State_0_sqmuxa, START_RNO_net_1, 
        N_79_i_0, NGRST_RNO_net_1, N_1369_i_0, Flag_Once_net_1, 
        Flag_Once_0_sqmuxa, \State[0]_net_1 , N_750_i_0, 
        \State[1]_net_1 , \State_ns[1] , \Byte_Count[0]_net_1 , 
        \Byte_Count_s[0] , N_753_i_0, \Byte_Count[1]_net_1 , 
        \Byte_Count_s[1] , \Byte_Count[2]_net_1 , \Byte_Count_s[2] , 
        \Byte_Count[3]_net_1 , \Byte_Count_s[3] , 
        \Byte_Count[4]_net_1 , \Byte_Count_s[4] , 
        \Byte_Count[5]_net_1 , \Byte_Count_s[5] , 
        \Byte_Count[6]_net_1 , \Byte_Count_s[6] , 
        \Byte_Count[7]_net_1 , \Byte_Count_s[7] , Byte_Count_cry_cy, 
        \State_RNIP3F3_Y[0] , \Byte_Count_cry[0] , \Byte_Count_cry[1] , 
        \Byte_Count_cry[2] , \Byte_Count_cry[3] , \Byte_Count_cry[4] , 
        \Byte_Count_cry[5] , \Byte_Count_cry[6] , N_1359, m11_i_0_a2_5, 
        m11_i_0_a2_4, N_1309;
    
    CFG4 #( .INIT(16'hCDCF) )  un1_State_0_sqmuxa_i_0_0_o2 (.A(ENCRC), 
        .B(\State[1]_net_1 ), .C(\State[0]_net_1 ), .D(TM_RSENC_0_RFS), 
        .Y(N_1309));
    ARI1 #( .INIT(20'h48800) )  \Byte_Count_RNO[7]  (.A(VCC_net_1), .B(
        \State_RNIP3F3_Y[0] ), .C(\Byte_Count[7]_net_1 ), .D(GND_net_1)
        , .FCI(\Byte_Count_cry[6] ), .S(\Byte_Count_s[7] ), .Y(), .FCO(
        ));
    SLE \DATAINP[3]  (.D(\Data_Buff[3]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(State_0_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RSControl_0_DATAINP[3]));
    CFG4 #( .INIT(16'h007F) )  \State_ns_1_0_.N_750_i  (.A(
        m11_i_0_a2_5), .B(m11_i_0_a2_4), .C(N_1359), .D(N_1309), .Y(
        N_750_i_0));
    CFG3 #( .INIT(8'h20) )  START_RNO (.A(ENCRC), .B(\State[0]_net_1 ), 
        .C(TM_RSENC_0_RFS), .Y(START_RNO_net_1));
    SLE \DATAINP[7]  (.D(\Data_Buff[7]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(State_0_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RSControl_0_DATAINP[7]));
    CFG3 #( .INIT(8'h18) )  \State_ns_1_0_.m14_0_0  (.A(TM_RSENC_0_RFD)
        , .B(\State[1]_net_1 ), .C(\State[0]_net_1 ), .Y(\State_ns[1] )
        );
    ARI1 #( .INIT(20'h48800) )  \Byte_Count_RNI31I22[4]  (.A(VCC_net_1)
        , .B(\State_RNIP3F3_Y[0] ), .C(\Byte_Count[4]_net_1 ), .D(
        GND_net_1), .FCI(\Byte_Count_cry[3] ), .S(\Byte_Count_s[4] ), 
        .Y(), .FCO(\Byte_Count_cry[4] ));
    CFG2 #( .INIT(4'h1) )  START_RNO_0 (.A(N_1359), .B(
        \State[1]_net_1 ), .Y(N_79_i_0));
    SLE \Data_Buff[1]  (.D(CPU_W_HDL_R_0_DataO[1]), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_75_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_Buff[1]_net_1 ));
    SLE \Byte_Count[4]  (.D(\Byte_Count_s[4] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_753_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Byte_Count[4]_net_1 ));
    SLE \DATAINP[0]  (.D(\Data_Buff[0]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(State_0_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RSControl_0_DATAINP[0]));
    VCC VCC (.Y(VCC_net_1));
    ARI1 #( .INIT(20'h46600) )  \State_RNIP3F3[0]  (.A(VCC_net_1), .B(
        \State[0]_net_1 ), .C(\State[1]_net_1 ), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(\State_RNIP3F3_Y[0] ), .FCO(
        Byte_Count_cry_cy));
    SLE \Data_Buff[2]  (.D(CPU_W_HDL_R_0_DataO[2]), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_75_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_Buff[2]_net_1 ));
    SLE Flag_Once (.D(VCC_net_1), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        Flag_Once_0_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Flag_Once_net_1));
    SLE \Byte_Count[7]  (.D(\Byte_Count_s[7] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_753_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Byte_Count[7]_net_1 ));
    SLE \Byte_Count[1]  (.D(\Byte_Count_s[1] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_753_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Byte_Count[1]_net_1 ));
    SLE \DATAINP[1]  (.D(\Data_Buff[1]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(State_0_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RSControl_0_DATAINP[1]));
    GND GND (.Y(GND_net_1));
    SLE \DATAINP[6]  (.D(\Data_Buff[6]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(State_0_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RSControl_0_DATAINP[6]));
    SLE \State[0]  (.D(N_750_i_0), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\State[0]_net_1 ));
    CFG2 #( .INIT(4'h4) )  NGRST_RNO (.A(\State[1]_net_1 ), .B(
        Flag_Once_net_1), .Y(NGRST_RNO_net_1));
    CFG2 #( .INIT(4'h2) )  un1_State_0_sqmuxa_i_0_0_a3 (.A(
        \State[0]_net_1 ), .B(TM_RSENC_0_RFD), .Y(N_1359));
    CFG4 #( .INIT(16'h0001) )  \State_ns_1_0_.m11_i_0_a2_5  (.A(
        \Byte_Count[3]_net_1 ), .B(\Byte_Count[2]_net_1 ), .C(
        \Byte_Count[1]_net_1 ), .D(\Byte_Count[0]_net_1 ), .Y(
        m11_i_0_a2_5));
    SLE \DATAINP[4]  (.D(\Data_Buff[4]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(State_0_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RSControl_0_DATAINP[4]));
    SLE \DATAINP[5]  (.D(\Data_Buff[5]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(State_0_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RSControl_0_DATAINP[5]));
    SLE \Data_Buff[3]  (.D(CPU_W_HDL_R_0_DataO[3]), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_75_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_Buff[3]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \Byte_Count_RNIV5UL1[3]  (.A(VCC_net_1)
        , .B(\State_RNIP3F3_Y[0] ), .C(\Byte_Count[3]_net_1 ), .D(
        GND_net_1), .FCI(\Byte_Count_cry[2] ), .S(\Byte_Count_s[3] ), 
        .Y(), .FCO(\Byte_Count_cry[3] ));
    CLKINT NGRST_RNIHQ59 (.A(NGRST_net_1), .Y(RSControl_0_NGRST));
    SLE \Data_Buff[6]  (.D(CPU_W_HDL_R_0_DataO[6]), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_75_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_Buff[6]_net_1 ));
    SLE \Data_Buff[7]  (.D(CPU_W_HDL_R_0_DataO[7]), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_75_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_Buff[7]_net_1 ));
    CFG2 #( .INIT(4'h9) )  \State_ns_1_0_.m12_0_x3_0_x2_i  (.A(
        \State[0]_net_1 ), .B(\State[1]_net_1 ), .Y(N_1369_i_0));
    CFG4 #( .INIT(16'h0080) )  \State_ns_1_0_.m11_i_0_a2_4  (.A(
        \Byte_Count[7]_net_1 ), .B(\Byte_Count[6]_net_1 ), .C(
        \Byte_Count[5]_net_1 ), .D(\Byte_Count[4]_net_1 ), .Y(
        m11_i_0_a2_4));
    SLE START (.D(START_RNO_net_1), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        N_79_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(RSControl_0_START));
    SLE \State[1]  (.D(\State_ns[1] ), .CLK(Bit_Count_16dec_i_1[3]), 
        .EN(VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\State[1]_net_1 ));
    SLE \DATAINP[2]  (.D(\Data_Buff[2]_net_1 ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(State_0_sqmuxa), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RSControl_0_DATAINP[2]));
    CFG3 #( .INIT(8'h20) )  State_0_sqmuxa_0_a3_0_a2_0_a2 (.A(
        TM_RSENC_0_RFD), .B(\State[1]_net_1 ), .C(\State[0]_net_1 ), 
        .Y(State_0_sqmuxa));
    SLE \Byte_Count[6]  (.D(\Byte_Count_s[6] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_753_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Byte_Count[6]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \Byte_Count_RNISBA91[2]  (.A(VCC_net_1)
        , .B(\State_RNIP3F3_Y[0] ), .C(\Byte_Count[2]_net_1 ), .D(
        GND_net_1), .FCI(\Byte_Count_cry[1] ), .S(\Byte_Count_s[2] ), 
        .Y(), .FCO(\Byte_Count_cry[2] ));
    SLE \Byte_Count[5]  (.D(\Byte_Count_s[5] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_753_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Byte_Count[5]_net_1 ));
    CFG4 #( .INIT(16'hFDFF) )  \State_RNI081H[0]  (.A(ENCRC), .B(
        \State[1]_net_1 ), .C(\State[0]_net_1 ), .D(TM_RSENC_0_RFS), 
        .Y(N_753_i_0));
    CFG3 #( .INIT(8'h01) )  Flag_Once_0_sqmuxa_0_a2_0_a2 (.A(
        \State[0]_net_1 ), .B(Flag_Once_net_1), .C(\State[1]_net_1 ), 
        .Y(Flag_Once_0_sqmuxa));
    ARI1 #( .INIT(20'h48800) )  \Byte_Count_RNI8T5F2[5]  (.A(VCC_net_1)
        , .B(\State_RNIP3F3_Y[0] ), .C(\Byte_Count[5]_net_1 ), .D(
        GND_net_1), .FCI(\Byte_Count_cry[4] ), .S(\Byte_Count_s[5] ), 
        .Y(), .FCO(\Byte_Count_cry[5] ));
    SLE \Byte_Count[3]  (.D(\Byte_Count_s[3] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_753_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Byte_Count[3]_net_1 ));
    SLE \Data_Buff[5]  (.D(CPU_W_HDL_R_0_DataO[5]), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_75_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_Buff[5]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \Byte_Count_RNIQIMS[1]  (.A(VCC_net_1), 
        .B(\State_RNIP3F3_Y[0] ), .C(\Byte_Count[1]_net_1 ), .D(
        GND_net_1), .FCI(\Byte_Count_cry[0] ), .S(\Byte_Count_s[1] ), 
        .Y(), .FCO(\Byte_Count_cry[1] ));
    SLE \Byte_Count[0]  (.D(\Byte_Count_s[0] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_753_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Byte_Count[0]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \Byte_Count_RNIEQPR2[6]  (.A(VCC_net_1)
        , .B(\State_RNIP3F3_Y[0] ), .C(\Byte_Count[6]_net_1 ), .D(
        GND_net_1), .FCI(\Byte_Count_cry[5] ), .S(\Byte_Count_s[6] ), 
        .Y(), .FCO(\Byte_Count_cry[6] ));
    SLE \Byte_Count[2]  (.D(\Byte_Count_s[2] ), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_753_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Byte_Count[2]_net_1 ));
    SLE NGRST (.D(NGRST_RNO_net_1), .CLK(Bit_Count_16dec_i_1[3]), .EN(
        N_1369_i_0), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(NGRST_net_1));
    SLE \Data_Buff[4]  (.D(CPU_W_HDL_R_0_DataO[4]), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_75_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_Buff[4]_net_1 ));
    ARI1 #( .INIT(20'h42800) )  \Byte_Count_RNIPQ2G[0]  (.A(VCC_net_1), 
        .B(\Byte_Count[0]_net_1 ), .C(\State[1]_net_1 ), .D(
        \State[0]_net_1 ), .FCI(Byte_Count_cry_cy), .S(
        \Byte_Count_s[0] ), .Y(), .FCO(\Byte_Count_cry[0] ));
    CFG2 #( .INIT(4'h1) )  un1_State_0_sqmuxa_i_0_0_o2_RNI74S8 (.A(
        N_1309), .B(N_1359), .Y(N_75_i_0));
    SLE \Data_Buff[0]  (.D(CPU_W_HDL_R_0_DataO[0]), .CLK(
        Bit_Count_16dec_i_1[3]), .EN(N_75_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Data_Buff[0]_net_1 ));
    
endmodule


module TC_Decode(
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       RX_GPIO1_c,
       C_1,
       FALG_FINISH_A_0,
       TC_Decode_0_IP_END_O,
       EnIP,
       RXRandomize_0_Block_ErrO,
       pending_0,
       ENCRC_0,
       RXRandomize_0_IP_END_O
    );
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  RX_GPIO1_c;
output C_1;
output FALG_FINISH_A_0;
output TC_Decode_0_IP_END_O;
output EnIP;
input  RXRandomize_0_Block_ErrO;
input  pending_0;
input  ENCRC_0;
input  RXRandomize_0_IP_END_O;

    wire \Bit_Count[4]_net_1 , VCC_net_1, N_801_i_0, Bit_Counte, 
        GND_net_1, \Bit_Count[1]_net_1 , N_804_i_0, 
        \Bit_Count[2]_net_1 , N_803_i_0, \Bit_Count[3]_net_1 , 
        N_802_i_0, \Bit_Count[0]_net_1 , N_815, 
        \HEAD_BUFFER[22]_net_1 , N_394, \Block_Count[0]_net_1 , 
        N_13_i_0, \Block_Count[1]_net_1 , N_788_i_0, 
        \Block_Count[2]_net_1 , N_787_i_0, \HEAD_BUFFER[7]_net_1 , 
        N_385, \HEAD_BUFFER[8]_net_1 , N_376, \HEAD_BUFFER[9]_net_1 , 
        HEAD_BUFFER_7_3_250_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[10]_net_1 , 
        HEAD_BUFFER_7_4_239_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[11]_net_1 , 
        HEAD_BUFFER_7_5_228_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[12]_net_1 , N_340, \HEAD_BUFFER[13]_net_1 , N_331, 
        \HEAD_BUFFER[14]_net_1 , N_322, \HEAD_BUFFER[15]_net_1 , N_313, 
        \HEAD_BUFFER[16]_net_1 , N_304, \HEAD_BUFFER[17]_net_1 , 
        HEAD_BUFFER_7_11_162_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[18]_net_1 , 
        HEAD_BUFFER_7_12_151_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[19]_net_1 , 
        HEAD_BUFFER_7_13_140_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[20]_net_1 , N_268, \HEAD_BUFFER[21]_net_1 , 
        HEAD_BUFFER_7_15_118_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[0]_net_1 , 
        HEAD_BUFFER_7_16_107_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[1]_net_1 , HEAD_BUFFER_7_17_96_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[2]_net_1 , HEAD_BUFFER_7_18_85_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[3]_net_1 , HEAD_BUFFER_7_19_74_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[4]_net_1 , HEAD_BUFFER_7_20_63_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[5]_net_1 , HEAD_BUFFER_7_21_52_a2_0_a4_0_a2_net_1, 
        \HEAD_BUFFER[6]_net_1 , HEAD_BUFFER_7_22_41_a2_0_a4_0_a2_net_1, 
        Head_error_net_1, N_800_i_0, Block_ErrO13_i_0, DataO_3, 
        IP_END_O_3_net_1, un1_Block_ErrO14_i_0, N_1110, N_1105, 
        Head_error_1_sqmuxa_i_0_a2_16_net_1, 
        Head_error_1_sqmuxa_i_0_a2_15_net_1, 
        Head_error_1_sqmuxa_i_0_a2_14_net_1, 
        Head_error_1_sqmuxa_i_0_a2_13_net_1, 
        Head_error_1_sqmuxa_i_0_a2_12_net_1, 
        Head_error_1_sqmuxa_i_0_a2_11_net_1, N_1102, 
        Head_error_1_sqmuxa_i_0_2_net_1, 
        Head_error_1_sqmuxa_i_0_a2_20_net_1;
    
    CFG4 #( .INIT(16'h00A6) )  \Block_Count_RNO[0]  (.A(
        \Block_Count[0]_net_1 ), .B(pending_0), .C(EnIP), .D(N_1110), 
        .Y(N_13_i_0));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_13_140_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[18]_net_1 ), .Y(
        HEAD_BUFFER_7_13_140_a2_0_a4_0_a2_net_1));
    SLE \HEAD_BUFFER[6]  (.D(HEAD_BUFFER_7_22_41_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[6]_net_1 ));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_18_85_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[1]_net_1 ), .Y(
        HEAD_BUFFER_7_18_85_a2_0_a4_0_a2_net_1));
    CFG4 #( .INIT(16'h0001) )  Head_error_1_sqmuxa_i_0_a2_16 (.A(
        \HEAD_BUFFER[14]_net_1 ), .B(\HEAD_BUFFER[5]_net_1 ), .C(
        \HEAD_BUFFER[2]_net_1 ), .D(\HEAD_BUFFER[0]_net_1 ), .Y(
        Head_error_1_sqmuxa_i_0_a2_16_net_1));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_6_217_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[11]_net_1 ), .Y(N_340));
    SLE IP_END_O (.D(IP_END_O_3_net_1), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(TC_Decode_0_IP_END_O));
    SLE Head_error (.D(N_800_i_0), .CLK(RX_GPIO1_c), .EN(VCC_net_1), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Head_error_net_1));
    SLE \Bit_Count[4]  (.D(N_801_i_0), .CLK(RX_GPIO1_c), .EN(
        Bit_Counte), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[4]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  Head_error_1_sqmuxa_i_0_a2_12 (.A(
        \HEAD_BUFFER[12]_net_1 ), .B(\HEAD_BUFFER[11]_net_1 ), .C(
        \HEAD_BUFFER[10]_net_1 ), .D(\HEAD_BUFFER[8]_net_1 ), .Y(
        Head_error_1_sqmuxa_i_0_a2_12_net_1));
    CFG3 #( .INIT(8'h01) )  Head_error_1_sqmuxa_i_0_a2_11 (.A(
        \HEAD_BUFFER[22]_net_1 ), .B(\HEAD_BUFFER[13]_net_1 ), .C(
        ENCRC_0), .Y(Head_error_1_sqmuxa_i_0_a2_11_net_1));
    SLE \HEAD_BUFFER[5]  (.D(HEAD_BUFFER_7_21_52_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[5]_net_1 ));
    SLE \HEAD_BUFFER[13]  (.D(N_331), .CLK(RX_GPIO1_c), .EN(Bit_Counte)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\HEAD_BUFFER[13]_net_1 ));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_1_272_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[6]_net_1 ), .Y(N_385));
    SLE \HEAD_BUFFER[15]  (.D(N_313), .CLK(RX_GPIO1_c), .EN(Bit_Counte)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\HEAD_BUFFER[15]_net_1 ));
    CFG2 #( .INIT(4'h2) )  Bit_Count_n0_i_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\Bit_Count[0]_net_1 ), .Y(N_815));
    SLE \Bit_Count[1]  (.D(N_804_i_0), .CLK(RX_GPIO1_c), .EN(
        Bit_Counte), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  Head_error_1_sqmuxa_i_0_o2 (.A(
        Block_ErrO13_i_0), .B(pending_0), .Y(un1_Block_ErrO14_i_0));
    CFG4 #( .INIT(16'h1333) )  Head_error_RNO (.A(
        Head_error_1_sqmuxa_i_0_a2_20_net_1), .B(
        Head_error_1_sqmuxa_i_0_2_net_1), .C(
        Head_error_1_sqmuxa_i_0_a2_16_net_1), .D(
        Head_error_1_sqmuxa_i_0_a2_15_net_1), .Y(N_800_i_0));
    SLE \HEAD_BUFFER[7]  (.D(N_385), .CLK(RX_GPIO1_c), .EN(Bit_Counte), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[7]_net_1 ));
    CFG2 #( .INIT(4'hE) )  Head_error_RNI4NE8 (.A(
        RXRandomize_0_Block_ErrO), .B(Head_error_net_1), .Y(
        Block_ErrO13_i_0));
    SLE \HEAD_BUFFER[1]  (.D(HEAD_BUFFER_7_17_96_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[1]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h4) )  IP_END_O_3 (.A(Block_ErrO13_i_0), .B(
        RXRandomize_0_IP_END_O), .Y(IP_END_O_3_net_1));
    SLE DataO (.D(DataO_3), .CLK(RX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        FALG_FINISH_A_0));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_5_228_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[10]_net_1 ), .Y(
        HEAD_BUFFER_7_5_228_a2_0_a4_0_a2_net_1));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_14_129_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[19]_net_1 ), .Y(N_268));
    CFG4 #( .INIT(16'h84C0) )  \Block_Count_RNO[2]  (.A(N_1105), .B(
        un1_Block_ErrO14_i_0), .C(\Block_Count[2]_net_1 ), .D(
        \Block_Count[1]_net_1 ), .Y(N_787_i_0));
    SLE \Block_Count[1]  (.D(N_788_i_0), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Block_Count[1]_net_1 ));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_7_206_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[12]_net_1 ), .Y(N_331));
    SLE \HEAD_BUFFER[3]  (.D(HEAD_BUFFER_7_19_74_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[3]_net_1 ));
    SLE Block_ErrO (.D(Block_ErrO13_i_0), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(C_1));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_2_261_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[7]_net_1 ), .Y(N_376));
    SLE \HEAD_BUFFER[0]  (.D(HEAD_BUFFER_7_16_107_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[0]_net_1 ));
    CFG4 #( .INIT(16'h84C0) )  \Bit_Count_RNO[4]  (.A(N_1102), .B(
        un1_Block_ErrO14_i_0), .C(\Bit_Count[4]_net_1 ), .D(
        \Bit_Count[3]_net_1 ), .Y(N_801_i_0));
    SLE \HEAD_BUFFER[2]  (.D(HEAD_BUFFER_7_18_85_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[2]_net_1 ));
    SLE \Block_Count[2]  (.D(N_787_i_0), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Block_Count[2]_net_1 ));
    SLE \Bit_Count[2]  (.D(N_803_i_0), .CLK(RX_GPIO1_c), .EN(
        Bit_Counte), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[2]_net_1 ));
    SLE \HEAD_BUFFER[4]  (.D(HEAD_BUFFER_7_20_63_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[4]_net_1 ));
    SLE \HEAD_BUFFER[14]  (.D(N_322), .CLK(RX_GPIO1_c), .EN(Bit_Counte)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\HEAD_BUFFER[14]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h0100) )  Head_error_1_sqmuxa_i_0_a2_13 (.A(
        \HEAD_BUFFER[19]_net_1 ), .B(\HEAD_BUFFER[18]_net_1 ), .C(
        \HEAD_BUFFER[9]_net_1 ), .D(\HEAD_BUFFER[4]_net_1 ), .Y(
        Head_error_1_sqmuxa_i_0_a2_13_net_1));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_9_184_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[14]_net_1 ), .Y(N_313));
    SLE \HEAD_BUFFER[19]  (.D(HEAD_BUFFER_7_13_140_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[19]_net_1 ));
    SLE En_DataO (.D(un1_Block_ErrO14_i_0), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(EnIP));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_22_41_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[5]_net_1 ), .Y(
        HEAD_BUFFER_7_22_41_a2_0_a4_0_a2_net_1));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_21_52_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[4]_net_1 ), .Y(
        HEAD_BUFFER_7_21_52_a2_0_a4_0_a2_net_1));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_10_173_a2_0_a4 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[15]_net_1 ), .Y(N_304));
    SLE \HEAD_BUFFER[20]  (.D(N_268), .CLK(RX_GPIO1_c), .EN(Bit_Counte)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\HEAD_BUFFER[20]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  Head_error_1_sqmuxa_i_0_a2_14 (.A(
        \HEAD_BUFFER[20]_net_1 ), .B(\HEAD_BUFFER[17]_net_1 ), .C(
        \HEAD_BUFFER[16]_net_1 ), .D(\HEAD_BUFFER[6]_net_1 ), .Y(
        Head_error_1_sqmuxa_i_0_a2_14_net_1));
    CFG2 #( .INIT(4'hB) )  \Block_Count_6_i_0_o2_1[0]  (.A(EnIP), .B(
        \Block_Count[0]_net_1 ), .Y(N_1105));
    SLE \HEAD_BUFFER[10]  (.D(HEAD_BUFFER_7_4_239_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[10]_net_1 ));
    SLE \HEAD_BUFFER[21]  (.D(HEAD_BUFFER_7_15_118_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[21]_net_1 ));
    CFG3 #( .INIT(8'h48) )  \Bit_Count_RNO[1]  (.A(
        \Bit_Count[0]_net_1 ), .B(un1_Block_ErrO14_i_0), .C(
        \Bit_Count[1]_net_1 ), .Y(N_804_i_0));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_17_96_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[0]_net_1 ), .Y(
        HEAD_BUFFER_7_17_96_a2_0_a4_0_a2_net_1));
    CFG4 #( .INIT(16'hCEEE) )  HEAD_BUFFER_1_sqmuxa_i_0_o2_0 (.A(
        pending_0), .B(N_1110), .C(\Bit_Count[4]_net_1 ), .D(
        \Bit_Count[3]_net_1 ), .Y(Bit_Counte));
    SLE \Bit_Count[0]  (.D(N_815), .CLK(RX_GPIO1_c), .EN(Bit_Counte), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Bit_Count[0]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  Head_error_1_sqmuxa_i_0_o2_0 (.A(
        \Bit_Count[2]_net_1 ), .B(\Bit_Count[1]_net_1 ), .C(
        \Bit_Count[0]_net_1 ), .Y(N_1102));
    SLE \HEAD_BUFFER[11]  (.D(HEAD_BUFFER_7_5_228_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[11]_net_1 ));
    SLE \HEAD_BUFFER[22]  (.D(N_394), .CLK(RX_GPIO1_c), .EN(Bit_Counte)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\HEAD_BUFFER[22]_net_1 ));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_8_195_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[13]_net_1 ), .Y(N_322));
    CFG4 #( .INIT(16'h48C0) )  \Bit_Count_RNO[2]  (.A(
        \Bit_Count[0]_net_1 ), .B(un1_Block_ErrO14_i_0), .C(
        \Bit_Count[2]_net_1 ), .D(\Bit_Count[1]_net_1 ), .Y(N_803_i_0));
    CFG4 #( .INIT(16'hFFBF) )  Head_error_1_sqmuxa_i_0_2 (.A(N_1102), 
        .B(un1_Block_ErrO14_i_0), .C(\Bit_Count[4]_net_1 ), .D(
        \Bit_Count[3]_net_1 ), .Y(Head_error_1_sqmuxa_i_0_2_net_1));
    SLE \HEAD_BUFFER[12]  (.D(N_340), .CLK(RX_GPIO1_c), .EN(Bit_Counte)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\HEAD_BUFFER[12]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  Head_error_1_sqmuxa_i_0_a2_20 (.A(
        Head_error_1_sqmuxa_i_0_a2_13_net_1), .B(
        Head_error_1_sqmuxa_i_0_a2_11_net_1), .C(
        Head_error_1_sqmuxa_i_0_a2_12_net_1), .D(
        Head_error_1_sqmuxa_i_0_a2_14_net_1), .Y(
        Head_error_1_sqmuxa_i_0_a2_20_net_1));
    CFG2 #( .INIT(4'h4) )  DataO_3_0_a2 (.A(Block_ErrO13_i_0), .B(
        ENCRC_0), .Y(DataO_3));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_16_107_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(ENCRC_0), .Y(
        HEAD_BUFFER_7_16_107_a2_0_a4_0_a2_net_1));
    SLE \HEAD_BUFFER[18]  (.D(HEAD_BUFFER_7_12_151_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[18]_net_1 ));
    CFG3 #( .INIT(8'h84) )  \Bit_Count_RNO[3]  (.A(N_1102), .B(
        un1_Block_ErrO14_i_0), .C(\Bit_Count[3]_net_1 ), .Y(N_802_i_0));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_3_250_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[8]_net_1 ), .Y(
        HEAD_BUFFER_7_3_250_a2_0_a4_0_a2_net_1));
    SLE \HEAD_BUFFER[9]  (.D(HEAD_BUFFER_7_3_250_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[9]_net_1 ));
    SLE \Block_Count[0]  (.D(N_13_i_0), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Block_Count[0]_net_1 ));
    CFG4 #( .INIT(16'hEEFE) )  HEAD_BUFFER_1_sqmuxa_i_0_o2_0_o2 (.A(
        RXRandomize_0_Block_ErrO), .B(Head_error_net_1), .C(
        \Block_Count[2]_net_1 ), .D(pending_0), .Y(N_1110));
    CFG4 #( .INIT(16'h00C6) )  \Block_Count_RNO[1]  (.A(pending_0), .B(
        \Block_Count[1]_net_1 ), .C(N_1105), .D(N_1110), .Y(N_788_i_0));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_11_162_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[16]_net_1 ), .Y(
        HEAD_BUFFER_7_11_162_a2_0_a4_0_a2_net_1));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_4_239_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[9]_net_1 ), .Y(
        HEAD_BUFFER_7_4_239_a2_0_a4_0_a2_net_1));
    SLE \HEAD_BUFFER[17]  (.D(HEAD_BUFFER_7_11_162_a2_0_a4_0_a2_net_1), 
        .CLK(RX_GPIO1_c), .EN(Bit_Counte), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[17]_net_1 ));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_15_118_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[20]_net_1 ), .Y(
        HEAD_BUFFER_7_15_118_a2_0_a4_0_a2_net_1));
    SLE \HEAD_BUFFER[16]  (.D(N_304), .CLK(RX_GPIO1_c), .EN(Bit_Counte)
        , .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\HEAD_BUFFER[16]_net_1 ));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_20_63_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[3]_net_1 ), .Y(
        HEAD_BUFFER_7_20_63_a2_0_a4_0_a2_net_1));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_19_74_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[2]_net_1 ), .Y(
        HEAD_BUFFER_7_19_74_a2_0_a4_0_a2_net_1));
    SLE \HEAD_BUFFER[8]  (.D(N_376), .CLK(RX_GPIO1_c), .EN(Bit_Counte), 
        .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \HEAD_BUFFER[8]_net_1 ));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_0_283_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[21]_net_1 ), .Y(N_394));
    CFG4 #( .INIT(16'h0001) )  Head_error_1_sqmuxa_i_0_a2_15 (.A(
        \HEAD_BUFFER[21]_net_1 ), .B(\HEAD_BUFFER[7]_net_1 ), .C(
        \HEAD_BUFFER[3]_net_1 ), .D(\HEAD_BUFFER[1]_net_1 ), .Y(
        Head_error_1_sqmuxa_i_0_a2_15_net_1));
    SLE \Bit_Count[3]  (.D(N_802_i_0), .CLK(RX_GPIO1_c), .EN(
        Bit_Counte), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\Bit_Count[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  HEAD_BUFFER_7_12_151_a2_0_a4_0_a2 (.A(
        un1_Block_ErrO14_i_0), .B(\HEAD_BUFFER[17]_net_1 ), .Y(
        HEAD_BUFFER_7_12_151_a2_0_a4_0_a2_net_1));
    
endmodule


module RXRandomize(
       test_4463andcpuopration_MSS_0_GPIO_1_M2F,
       RX_GPIO1_c,
       ENCRC_0,
       pending_0,
       RXRandomize_0_Block_ErrO,
       CLTU_0_Block_ErrO,
       RXRandomize_0_IP_END_O,
       CLTU_0_IP_END,
       ENASM_0,
       A_1
    );
input  test_4463andcpuopration_MSS_0_GPIO_1_M2F;
input  RX_GPIO1_c;
output ENCRC_0;
output pending_0;
output RXRandomize_0_Block_ErrO;
input  CLTU_0_Block_ErrO;
output RXRandomize_0_IP_END_O;
input  CLTU_0_IP_END;
input  ENASM_0;
input  A_1;

    wire \Ran_SR[4]_net_1 , GND_net_1, N_238_i_0, 
        un1_Ran_SR30_2_i_0_net_1, VCC_net_1, \Ran_SR[5]_net_1 , 
        N_229_i_0, \Ran_SR[6]_net_1 , N_220_i_0, \Ran_SR[7]_net_1 , 
        N_766_i_0, \Start_Buff[5]_net_1 , \Start_Buff_5[5] , 
        un1_Block_ErrI_3_i_0, \Start_Buff[6]_net_1 , \Start_Buff_5[6] , 
        \Start_Buff[7]_net_1 , \Start_Buff_5[7] , 
        \Start_Buff[8]_net_1 , \Start_Buff_5[8] , 
        \Start_Buff[9]_net_1 , \Start_Buff_5[9] , 
        \Start_Buff[10]_net_1 , \Start_Buff_5[10] , 
        \Start_Buff[11]_net_1 , \Start_Buff_5[11] , 
        \Start_Buff[12]_net_1 , \Start_Buff_5[12] , 
        \Start_Buff[13]_net_1 , \Start_Buff_5[13] , 
        \Start_Buff[14]_net_1 , \Start_Buff_5[14] , 
        \Start_Buff[15]_net_1 , \Start_Buff_5[15] , \Ran_SR[0]_net_1 , 
        N_184_i_0, \Ran_SR[1]_net_1 , N_175_i_0, \Ran_SR[2]_net_1 , 
        N_166_i_0, \Ran_SR[3]_net_1 , N_157_i_0, \Start_Buff[0]_net_1 , 
        \Start_Buff_5[0] , \Start_Buff[1]_net_1 , \Start_Buff_5[1] , 
        \Start_Buff[2]_net_1 , \Start_Buff_5[2] , 
        \Start_Buff[3]_net_1 , \Start_Buff_5[3] , 
        \Start_Buff[4]_net_1 , \Start_Buff_5[4] , N_145_i_0, 
        un1_Ran_SR30_i_0_net_1, N_760_i_0, Flag_once_net_1, N_764_i_0, 
        N_17, Ran_SR30, N_771, N_763, un1_Block_ErrI_3_0_a2_11_net_1, 
        un1_Block_ErrI_3_0_a2_10_net_1, un1_Block_ErrI_3_0_a2_9_net_1, 
        un1_Block_ErrI_3_0_a2_8_net_1, Ran_SR_11_2_110_x2_3_net_1, 
        N_786;
    
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[3]  (.A(
        \Start_Buff[2]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[3] ));
    SLE \Start_Buff[2]  (.D(\Start_Buff_5[2] ), .CLK(RX_GPIO1_c), .EN(
        un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[10]  (.A(
        \Start_Buff[9]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[10] ));
    SLE \Start_Buff[9]  (.D(\Start_Buff_5[9] ), .CLK(RX_GPIO1_c), .EN(
        un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[9]_net_1 ));
    SLE EnO (.D(N_760_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_Ran_SR30_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(pending_0)
        );
    SLE IP_END_O (.D(Ran_SR30), .CLK(RX_GPIO1_c), .EN(VCC_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RXRandomize_0_IP_END_O));
    SLE \Ran_SR[4]  (.D(N_238_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_Ran_SR30_2_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Ran_SR[4]_net_1 ));
    SLE \Start_Buff[4]  (.D(\Start_Buff_5[4] ), .CLK(RX_GPIO1_c), .EN(
        un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[4]_net_1 ));
    CFG2 #( .INIT(4'h1) )  Flag_once_RNO (.A(CLTU_0_Block_ErrO), .B(
        CLTU_0_IP_END), .Y(N_764_i_0));
    SLE \Start_Buff[3]  (.D(\Start_Buff_5[3] ), .CLK(RX_GPIO1_c), .EN(
        un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[3]_net_1 ));
    CFG4 #( .INIT(16'hFF40) )  un1_Ran_SR30_i_0 (.A(CLTU_0_IP_END), .B(
        Flag_once_net_1), .C(N_786), .D(CLTU_0_Block_ErrO), .Y(
        un1_Ran_SR30_i_0_net_1));
    CFG2 #( .INIT(4'hD) )  \Ran_SR_RNO[3]  (.A(N_771), .B(
        \Ran_SR[4]_net_1 ), .Y(N_157_i_0));
    CFG4 #( .INIT(16'hFFBA) )  un1_Block_ErrI_5_i_0 (.A(CLTU_0_IP_END), 
        .B(Flag_once_net_1), .C(N_786), .D(CLTU_0_Block_ErrO), .Y(N_17)
        );
    SLE \Ran_SR[3]  (.D(N_157_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_Ran_SR30_2_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Ran_SR[3]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  un1_Block_ErrI_3_0_a2_9 (.A(
        \Start_Buff[12]_net_1 ), .B(\Start_Buff[6]_net_1 ), .C(
        \Start_Buff[5]_net_1 ), .D(\Start_Buff[2]_net_1 ), .Y(
        un1_Block_ErrI_3_0_a2_9_net_1));
    SLE \Start_Buff[6]  (.D(\Start_Buff_5[6] ), .CLK(RX_GPIO1_c), .EN(
        un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[6]_net_1 ));
    SLE \Start_Buff[15]  (.D(\Start_Buff_5[15] ), .CLK(RX_GPIO1_c), 
        .EN(un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[15]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[11]  (.A(
        \Start_Buff[10]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[11] ));
    VCC VCC (.Y(VCC_net_1));
    SLE DataO (.D(N_145_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_Ran_SR30_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(ENCRC_0));
    SLE \Start_Buff[8]  (.D(\Start_Buff_5[8] ), .CLK(RX_GPIO1_c), .EN(
        un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[8]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  un1_Block_ErrI_3_0_a2_8 (.A(
        \Start_Buff[15]_net_1 ), .B(\Start_Buff[3]_net_1 ), .C(
        \Start_Buff[1]_net_1 ), .D(\Start_Buff[0]_net_1 ), .Y(
        un1_Block_ErrI_3_0_a2_8_net_1));
    SLE \Ran_SR[5]  (.D(N_229_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_Ran_SR30_2_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Ran_SR[5]_net_1 ));
    SLE Block_ErrO (.D(CLTU_0_Block_ErrO), .CLK(RX_GPIO1_c), .EN(
        VCC_net_1), .ALn(test_4463andcpuopration_MSS_0_GPIO_1_M2F), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(RXRandomize_0_Block_ErrO));
    SLE \Ran_SR[7]  (.D(N_766_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_Ran_SR30_2_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Ran_SR[7]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[4]  (.A(
        \Start_Buff[3]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[4] ));
    SLE \Start_Buff[1]  (.D(\Start_Buff_5[1] ), .CLK(RX_GPIO1_c), .EN(
        un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[1]_net_1 ));
    SLE Flag_once (.D(N_764_i_0), .CLK(RX_GPIO1_c), .EN(N_17), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Flag_once_net_1));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[2]  (.A(
        \Start_Buff[1]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[2] ));
    CFG4 #( .INIT(16'h0080) )  un1_Block_ErrI_3_0_a2_10 (.A(
        \Start_Buff[14]_net_1 ), .B(\Start_Buff[13]_net_1 ), .C(
        \Start_Buff[11]_net_1 ), .D(\Start_Buff[10]_net_1 ), .Y(
        un1_Block_ErrI_3_0_a2_10_net_1));
    SLE \Start_Buff[7]  (.D(\Start_Buff_5[7] ), .CLK(RX_GPIO1_c), .EN(
        un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[7]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \Start_Buff[14]  (.D(\Start_Buff_5[14] ), .CLK(RX_GPIO1_c), 
        .EN(un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[14]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \Ran_SR_RNO[6]  (.A(N_771), .B(
        \Ran_SR[7]_net_1 ), .Y(N_220_i_0));
    SLE \Ran_SR[6]  (.D(N_220_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_Ran_SR30_2_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Ran_SR[6]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[5]  (.A(
        \Start_Buff[4]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[5] ));
    CFG2 #( .INIT(4'h4) )  EnO_RNO (.A(CLTU_0_Block_ErrO), .B(ENASM_0), 
        .Y(N_760_i_0));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[14]  (.A(
        \Start_Buff[13]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[14] ));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[8]  (.A(
        \Start_Buff[7]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[8] ));
    CFG2 #( .INIT(4'hD) )  \Ran_SR_RNO[5]  (.A(N_771), .B(
        \Ran_SR[6]_net_1 ), .Y(N_229_i_0));
    CFG2 #( .INIT(4'hD) )  un1_Ran_SR30_2_i_o2 (.A(Flag_once_net_1), 
        .B(ENASM_0), .Y(N_763));
    CFG2 #( .INIT(4'hD) )  \Ran_SR_RNO[2]  (.A(N_771), .B(
        \Ran_SR[3]_net_1 ), .Y(N_166_i_0));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[7]  (.A(
        \Start_Buff[6]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[7] ));
    SLE \Start_Buff[11]  (.D(\Start_Buff_5[11] ), .CLK(RX_GPIO1_c), 
        .EN(un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[11]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[13]  (.A(
        \Start_Buff[12]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[13] ));
    CFG2 #( .INIT(4'hD) )  \Ran_SR_RNO[4]  (.A(N_771), .B(
        \Ran_SR[5]_net_1 ), .Y(N_238_i_0));
    CFG2 #( .INIT(4'hD) )  \Ran_SR_RNO[0]  (.A(N_771), .B(
        \Ran_SR[1]_net_1 ), .Y(N_184_i_0));
    CFG3 #( .INIT(8'hFB) )  un1_Block_ErrI_3_0_a2_RNID8511 (.A(
        CLTU_0_Block_ErrO), .B(N_786), .C(CLTU_0_IP_END), .Y(
        un1_Block_ErrI_3_i_0));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[6]  (.A(
        \Start_Buff[5]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[6] ));
    CFG4 #( .INIT(16'hB77B) )  \Ran_SR_RNO[7]  (.A(
        Ran_SR_11_2_110_x2_3_net_1), .B(N_771), .C(\Ran_SR[3]_net_1 ), 
        .D(\Ran_SR[2]_net_1 ), .Y(N_766_i_0));
    CFG2 #( .INIT(4'h4) )  Ran_SR30_0_a3 (.A(CLTU_0_Block_ErrO), .B(
        CLTU_0_IP_END), .Y(Ran_SR30));
    SLE \Start_Buff[5]  (.D(\Start_Buff_5[5] ), .CLK(RX_GPIO1_c), .EN(
        un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[5]_net_1 ));
    SLE \Start_Buff[0]  (.D(\Start_Buff_5[0] ), .CLK(RX_GPIO1_c), .EN(
        un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[0]_net_1 ));
    CFG4 #( .INIT(16'h0220) )  DataO_RNO (.A(ENASM_0), .B(
        CLTU_0_Block_ErrO), .C(\Ran_SR[0]_net_1 ), .D(A_1), .Y(
        N_145_i_0));
    CFG4 #( .INIT(16'h8000) )  un1_Block_ErrI_3_0_a2 (.A(
        un1_Block_ErrI_3_0_a2_11_net_1), .B(
        un1_Block_ErrI_3_0_a2_10_net_1), .C(
        un1_Block_ErrI_3_0_a2_9_net_1), .D(
        un1_Block_ErrI_3_0_a2_8_net_1), .Y(N_786));
    CFG3 #( .INIT(8'h04) )  \Start_Buff_5_0_a3[0]  (.A(
        CLTU_0_Block_ErrO), .B(A_1), .C(CLTU_0_IP_END), .Y(
        \Start_Buff_5[0] ));
    CFG2 #( .INIT(4'h4) )  Ran_SR_11_0_159_i_a2_0_a2 (.A(
        CLTU_0_Block_ErrO), .B(Flag_once_net_1), .Y(N_771));
    SLE \Ran_SR[2]  (.D(N_166_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_Ran_SR30_2_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Ran_SR[2]_net_1 ));
    CFG4 #( .INIT(16'h6996) )  Ran_SR_11_2_110_x2_3 (.A(
        \Ran_SR[6]_net_1 ), .B(\Ran_SR[4]_net_1 ), .C(
        \Ran_SR[1]_net_1 ), .D(\Ran_SR[0]_net_1 ), .Y(
        Ran_SR_11_2_110_x2_3_net_1));
    SLE \Ran_SR[1]  (.D(N_175_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_Ran_SR30_2_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Ran_SR[1]_net_1 ));
    SLE \Start_Buff[12]  (.D(\Start_Buff_5[12] ), .CLK(RX_GPIO1_c), 
        .EN(un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[12]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  un1_Block_ErrI_3_0_a2_11 (.A(
        \Start_Buff[9]_net_1 ), .B(\Start_Buff[8]_net_1 ), .C(
        \Start_Buff[7]_net_1 ), .D(\Start_Buff[4]_net_1 ), .Y(
        un1_Block_ErrI_3_0_a2_11_net_1));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[9]  (.A(
        \Start_Buff[8]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[9] ));
    SLE \Start_Buff[10]  (.D(\Start_Buff_5[10] ), .CLK(RX_GPIO1_c), 
        .EN(un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[10]_net_1 ));
    SLE \Start_Buff[13]  (.D(\Start_Buff_5[13] ), .CLK(RX_GPIO1_c), 
        .EN(un1_Block_ErrI_3_i_0), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Start_Buff[13]_net_1 ));
    CFG2 #( .INIT(4'hD) )  \Ran_SR_RNO[1]  (.A(N_771), .B(
        \Ran_SR[2]_net_1 ), .Y(N_175_i_0));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[15]  (.A(
        \Start_Buff[14]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[15] ));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[12]  (.A(
        \Start_Buff[11]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[12] ));
    CFG4 #( .INIT(16'hAEAA) )  un1_Ran_SR30_2_i_0 (.A(
        CLTU_0_Block_ErrO), .B(N_786), .C(CLTU_0_IP_END), .D(N_763), 
        .Y(un1_Ran_SR30_2_i_0_net_1));
    CFG3 #( .INIT(8'h02) )  \Start_Buff_5_0_a3[1]  (.A(
        \Start_Buff[0]_net_1 ), .B(CLTU_0_IP_END), .C(
        CLTU_0_Block_ErrO), .Y(\Start_Buff_5[1] ));
    SLE \Ran_SR[0]  (.D(N_184_i_0), .CLK(RX_GPIO1_c), .EN(
        un1_Ran_SR30_2_i_0_net_1), .ALn(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \Ran_SR[0]_net_1 ));
    
endmodule


module test_4463andcpuopration(
       ADC_INT,
       BOARD_NO,
       CAN1_TX,
       CCA_NIRQ,
       DEVRST_N,
       L4V_PG,
       RXD4,
       RX_GPIO0,
       RX_GPIO1,
       SPI_MISO,
       TX_GPIO1,
       XTL,
       \A3.3V_EN ,
       ADC_CS,
       ADC_CSTART,
       ADC_FS,
       ADC_PWDN,
       ANT_SW1,
       ANT_SW2,
       CAN1_RS,
       CAN1_RX,
       CAN2_RS,
       L3V3_EN1,
       L3V3_EN2,
       L4463_RX_CS,
       L4463_TX_CS,
       L4V_EN,
       PA4V_ON,
       RX_SDN,
       SPI_CLK,
       SPI_FRAM_CS,
       SPI_MOSI,
       SW,
       TXD4,
       TX_GPIO0,
       TX_SDN
    );
input  ADC_INT;
input  BOARD_NO;
input  CAN1_TX;
input  CCA_NIRQ;
input  DEVRST_N;
input  L4V_PG;
input  RXD4;
input  RX_GPIO0;
input  RX_GPIO1;
input  SPI_MISO;
input  TX_GPIO1;
input  XTL;
output \A3.3V_EN ;
output ADC_CS;
output ADC_CSTART;
output ADC_FS;
output ADC_PWDN;
output ANT_SW1;
output ANT_SW2;
output CAN1_RS;
output CAN1_RX;
output CAN2_RS;
output L3V3_EN1;
output L3V3_EN2;
output L4463_RX_CS;
output L4463_TX_CS;
output L4V_EN;
output PA4V_ON;
output RX_SDN;
output SPI_CLK;
output SPI_FRAM_CS;
output SPI_MOSI;
output SW;
output TXD4;
output TX_GPIO0;
output TX_SDN;

    wire GND_net_1, VCC_net_1, P_CLK, 
        test_4463andcpuopration_MSS_0_GPIO_1_M2F, ENASM, ASM_OUT, 
        pending, A_1, ENASM_0, CLTU_0_Block_ErrO, CLTU_0_IP_END, 
        \CLTU_0_TC_Error_Counter[0] , CLTU_0_Flag_RX_ing, 
        Switch_0_EnOut, c_in, \CoreAPB3_0_APBmslave3_PADDR[0] , 
        \CoreAPB3_0_APBmslave3_PADDR[1] , 
        \CoreAPB3_0_APBmslave3_PADDR[9] , 
        \CoreAPB3_0_APBmslave3_PADDR[10] , 
        \CoreAPB3_0_APBmslave3_PADDR[11] , 
        \CoreAPB3_0_APBmslave3_PADDR[12] , 
        \CoreAPB3_0_APBmslave3_PADDR[13] , 
        \CoreAPB3_0_APBmslave3_PADDR[14] , 
        \CoreAPB3_0_APBmslave3_PADDR[15] , 
        \CoreAPB3_0_APBmslave3_PADDR[16] , 
        \CoreAPB3_0_APBmslave3_PADDR[17] , 
        \CoreAPB3_0_APBmslave3_PADDR[18] , 
        \CoreAPB3_0_APBmslave3_PADDR[19] , 
        \CoreAPB3_0_APBmslave3_PADDR[20] , 
        \CoreAPB3_0_APBmslave3_PADDR[21] , 
        \CoreAPB3_0_APBmslave3_PADDR[22] , 
        \CoreAPB3_0_APBmslave3_PADDR[23] , 
        \CoreAPB3_0_APBmslave3_PADDR[24] , 
        \CoreAPB3_0_APBmslave3_PADDR[25] , 
        \CoreAPB3_0_APBmslave3_PADDR[26] , 
        \CoreAPB3_0_APBmslave3_PADDR[27] , 
        \CoreAPB3_0_APBmslave3_PADDR[28] , 
        \CoreAPB3_0_APBmslave3_PADDR[29] , 
        \CoreAPB3_0_APBmslave3_PADDR[30] , 
        \CoreAPB3_0_APBmslave3_PADDR[31] , 
        CoreAPB3_0_APBmslave3_PWRITE, CoreAPB3_0_APBmslave3_PENABLE, 
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx, 
        \CoreAPB3_0_APBmslave3_PWDATA[0] , 
        \CoreAPB3_0_APBmslave3_PWDATA[1] , 
        \CoreAPB3_0_APBmslave3_PWDATA[2] , 
        \CoreAPB3_0_APBmslave3_PWDATA[3] , 
        \CoreAPB3_0_APBmslave3_PWDATA[4] , 
        \CoreAPB3_0_APBmslave3_PWDATA[5] , 
        \CoreAPB3_0_APBmslave3_PWDATA[6] , 
        \CoreAPB3_0_APBmslave3_PWDATA[7] , 
        \CoreAPB3_0_APBmslave3_PWDATA[8] , 
        \CoreAPB3_0_APBmslave3_PWDATA[9] , 
        \CoreAPB3_0_APBmslave3_PWDATA[10] , 
        \CoreAPB3_0_APBmslave3_PWDATA[11] , 
        \CoreAPB3_0_APBmslave3_PWDATA[12] , 
        \CoreAPB3_0_APBmslave3_PWDATA[13] , 
        \CoreAPB3_0_APBmslave3_PWDATA[14] , 
        \CoreAPB3_0_APBmslave3_PWDATA[15] , 
        \CoreAPB3_0_APBmslave3_PWDATA[16] , 
        \CoreAPB3_0_APBmslave3_PWDATA[17] , 
        \CoreAPB3_0_APBmslave3_PWDATA[18] , 
        \CoreAPB3_0_APBmslave3_PWDATA[19] , 
        \CoreAPB3_0_APBmslave3_PWDATA[20] , 
        \CoreAPB3_0_APBmslave3_PWDATA[21] , 
        \CoreAPB3_0_APBmslave3_PWDATA[22] , 
        \CoreAPB3_0_APBmslave3_PWDATA[23] , 
        \CoreAPB3_0_APBmslave3_PWDATA[24] , 
        \CoreAPB3_0_APBmslave3_PWDATA[25] , 
        \CoreAPB3_0_APBmslave3_PWDATA[26] , 
        \CoreAPB3_0_APBmslave3_PWDATA[27] , 
        \CoreAPB3_0_APBmslave3_PWDATA[28] , 
        \CoreAPB3_0_APBmslave3_PWDATA[29] , 
        \CoreAPB3_0_APBmslave3_PWDATA[30] , 
        \CoreAPB3_0_APBmslave3_PWDATA[31] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[0] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[16] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[17] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[18] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[19] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[20] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[21] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[22] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[23] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[24] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[25] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[26] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[27] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[28] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[29] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[30] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[31] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        \CoreAPB3_0_APBmslave3_PRDATA[8] , 
        \CoreAPB3_0_APBmslave3_PRDATA[9] , 
        \CoreAPB3_0_APBmslave3_PRDATA[10] , 
        \CoreAPB3_0_APBmslave3_PRDATA[11] , 
        \CoreAPB3_0_APBmslave3_PRDATA[12] , 
        \CoreAPB3_0_APBmslave3_PRDATA[13] , 
        \CoreAPB3_0_APBmslave3_PRDATA[14] , 
        \CoreAPB3_0_APBmslave3_PRDATA[15] , 
        \CoreAPB3_0_APBmslave3_PRDATA[16] , 
        \CoreAPB3_0_APBmslave3_PRDATA[17] , 
        \CoreAPB3_0_APBmslave3_PRDATA[18] , 
        \CoreAPB3_0_APBmslave3_PRDATA[19] , 
        \CoreAPB3_0_APBmslave3_PRDATA[20] , 
        \CoreAPB3_0_APBmslave3_PRDATA[21] , 
        \CoreAPB3_0_APBmslave3_PRDATA[22] , 
        \CoreAPB3_0_APBmslave3_PRDATA[23] , 
        \CoreAPB3_0_APBmslave3_PRDATA[24] , 
        \CoreAPB3_0_APBmslave3_PRDATA[25] , 
        \CoreAPB3_0_APBmslave3_PRDATA[26] , 
        \CoreAPB3_0_APBmslave3_PRDATA[27] , 
        \CoreAPB3_0_APBmslave3_PRDATA[28] , 
        \CoreAPB3_0_APBmslave3_PRDATA[29] , 
        \CoreAPB3_0_APBmslave3_PRDATA[30] , 
        \CoreAPB3_0_APBmslave3_PRDATA[31] , 
        CoreAPB3_0_APBmslave3_PREADY, OSC_0_XTLOSC_O2F, 
        \CPU_W_HDL_R_0_DataO[0] , \CPU_W_HDL_R_0_DataO[1] , 
        \CPU_W_HDL_R_0_DataO[2] , \CPU_W_HDL_R_0_DataO[3] , 
        \CPU_W_HDL_R_0_DataO[4] , \CPU_W_HDL_R_0_DataO[5] , 
        \CPU_W_HDL_R_0_DataO[6] , \CPU_W_HDL_R_0_DataO[7] , 
        Glue_Logic_0_USER_WEN_TRP1, \Glue_Logic_0_MSG_TRP1[0] , 
        \Glue_Logic_0_MSG_TRP1[1] , \Glue_Logic_0_MSG_TRP1[2] , 
        \Glue_Logic_0_MSG_TRP1[3] , \Glue_Logic_0_MSG_TRP1[4] , 
        \Glue_Logic_0_MSG_TRP1[5] , \Glue_Logic_0_MSG_TRP1[6] , 
        \Glue_Logic_0_MSG_TRP1[7] , \Glue_Logic_0_MSG_WA_TRP1[0] , 
        \Glue_Logic_0_MSG_WA_TRP1[1] , \Glue_Logic_0_MSG_WA_TRP1[2] , 
        \Glue_Logic_0_MSG_WA_TRP1[3] , \Glue_Logic_0_MSG_WA_TRP1[4] , 
        \Glue_Logic_0_MSG_WA_TRP1[5] , \Glue_Logic_0_MSG_WA_TRP1[6] , 
        \Glue_Logic_0_MSG_WA_TRP1[7] , \Glue_Logic_0_MSG_WA_TRP1[8] , 
        \Glue_Logic_0_MSG_WA_TRP1[9] , CPU_W_HDL_R_0_USER_REN_TRP1, 
        \CPU_W_HDL_R_0_USER_RA_TRP1[0] , 
        \CPU_W_HDL_R_0_USER_RA_TRP1[1] , 
        \CPU_W_HDL_R_0_USER_RA_TRP1[2] , 
        \CPU_W_HDL_R_0_USER_RA_TRP1[3] , 
        \CPU_W_HDL_R_0_USER_RA_TRP1[4] , 
        \CPU_W_HDL_R_0_USER_RA_TRP1[5] , 
        \CPU_W_HDL_R_0_USER_RA_TRP1[6] , 
        \CPU_W_HDL_R_0_USER_RA_TRP1[7] , 
        \CPU_W_HDL_R_0_USER_RA_TRP1[9] , 
        HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1, 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[0] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[1] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[2] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[3] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[4] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[5] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[6] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[7] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[8] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[9] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[10] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[11] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[12] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[13] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[14] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[15] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[16] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[17] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[18] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[19] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[20] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[21] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[22] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[23] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[24] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[25] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[26] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[27] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[28] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[29] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[30] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[31] , 
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0] , 
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[1] , 
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[2] , 
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[3] , 
        Glue_Logic_0_USER_REN_TRP1, \Glue_Logic_0_USER_RA_TRP1_1[0] , 
        \Glue_Logic_0_USER_RA_TRP1_1[1] , 
        \Glue_Logic_0_USER_RA_TRP1_1[2] , 
        \Glue_Logic_0_USER_RA_TRP1_1[3] , TXD4_net_0, 
        Glue_Logic_0_Flag_B_Tx, En_read_buff, 
        CPU_W_HDL_R_0_Flag_A_Tx_Finish, CPU_W_HDL_R_0_Flag_B_Tx_Finish, 
        ENCRC, \Glue_Logic_0_Flag_Int_0[0] , 
        HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish, 
        HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish, Flag_RX, 
        Glue_Logic_0_Flag_B_Rx, FALG_FINISH_A_0, EnIP, C_1, 
        TC_Decode_0_IP_END_O, 
        test_4463andcpuopration_MSS_0_GPIO_15_M2F, TM_RSENC_0_RDY, 
        \TM_RSENC_0_CODEOUTP[0] , \TM_RSENC_0_CODEOUTP[1] , 
        \TM_RSENC_0_CODEOUTP[2] , \TM_RSENC_0_CODEOUTP[3] , 
        \TM_RSENC_0_CODEOUTP[4] , \TM_RSENC_0_CODEOUTP[5] , 
        \TM_RSENC_0_CODEOUTP[6] , \TM_RSENC_0_CODEOUTP[7] , P_OUT, 
        S_OUT_0, TM_RSENC_0_RFD, TM_RSENC_0_RFS, RSControl_0_NGRST, 
        RSControl_0_START, \RSControl_0_DATAINP[0] , 
        \RSControl_0_DATAINP[1] , \RSControl_0_DATAINP[2] , 
        \RSControl_0_DATAINP[3] , \RSControl_0_DATAINP[4] , 
        \RSControl_0_DATAINP[5] , \RSControl_0_DATAINP[6] , 
        \RSControl_0_DATAINP[7] , ENCRC_0, pending_0, 
        RXRandomize_0_Block_ErrO, RXRandomize_0_IP_END_O, 
        SYSRESET_0_POWER_ON_RESET_N, \Randomizer_0.pn_reg[0] , 
        \Convolutional_Encoder_0.shift1_reg[4] , 
        \Convolutional_Encoder_0.shift1_reg[0] , 
        \ASM_Generato_0.stream[0] , ADC_INT_c, BOARD_NO_c, CAN1_TX_c, 
        CCA_NIRQ_c, L4V_PG_c, RXD4_c, RX_GPIO0_c, RX_GPIO1_c, 
        SPI_MISO_c, TX_GPIO1_c, \A3.3V_EN_c , ADC_CS_c, ADC_CSTART_c, 
        ADC_FS_c, ADC_PWDN_c, ANT_SW1_c, ANT_SW2_c, CAN1_RX_c, 
        L3V3_EN1_c, L3V3_EN2_c, L4463_RX_CS_c, L4463_TX_CS_c, L4V_EN_c, 
        PA4V_ON_c, RX_SDN_c, SPI_CLK_c, SPI_FRAM_CS_c, SPI_MOSI_c, 
        SW_c, TXD4_c, TX_GPIO0_c, TX_SDN_c, \COREEDAC_1_DATA_OUT[16] , 
        \COREEDAC_1_DATA_OUT[2] , \COREEDAC_1_DATA_OUT[4] , 
        \COREEDAC_1_DATA_OUT[10] , \COREEDAC_1_DATA_OUT[11] , 
        \COREEDAC_1_DATA_OUT[13] , \COREEDAC_1_DATA_OUT[28] , 
        \COREEDAC_1_DATA_OUT[24] , \COREEDAC_1_DATA_OUT[15] , 
        \COREEDAC_1_DATA_OUT[20] , \COREEDAC_1_DATA_OUT[12] , 
        \COREEDAC_1_DATA_OUT[1] , \COREEDAC_1_DATA_OUT[6] , 
        \COREEDAC_1_DATA_OUT[3] , \COREEDAC_1_DATA_OUT[25] , 
        \CoreAPB3_0.iPSELS_raw23 , \COREEDAC_1_DATA_OUT[29] , 
        \COREEDAC_1_DATA_OUT[26] , \COREEDAC_1_DATA_OUT[19] , 
        \COREEDAC_1_DATA_OUT[14] , \COREEDAC_1_DATA_OUT[7] , 
        \COREEDAC_1_DATA_OUT[8] , \COREEDAC_1_DATA_OUT[18] , 
        \COREEDAC_1_DATA_OUT[31] , \COREEDAC_1_DATA_OUT[22] , 
        \COREEDAC_1_DATA_OUT[21] , \COREEDAC_1_DATA_OUT[9] , 
        \COREEDAC_1_DATA_OUT[0] , \COREEDAC_1_DATA_OUT[30] , 
        \COREEDAC_1_DATA_OUT[5] , \COREEDAC_1_DATA_OUT[17] , 
        \COREEDAC_1_DATA_OUT[27] , \COREEDAC_1_DATA_OUT[23] , 
        \CoreAPB3_0_APBmslave3_PADDR[2] , 
        \CoreAPB3_0_APBmslave3_PADDR[3] , 
        \CoreAPB3_0_APBmslave3_PADDR[4] , 
        \CoreAPB3_0_APBmslave3_PADDR[5] , 
        \CoreAPB3_0_APBmslave3_PADDR[6] , 
        \CoreAPB3_0_APBmslave3_PADDR[7] , 
        \CoreAPB3_0_APBmslave3_PADDR[8] , 
        \Convolutional_Encoder_0.Convolutional_Encoder_out_1_0 , 
        \CLTU_0_TC_Packet_Counter[0] , \CLTU_0_TC_Packet_Counter[1] , 
        \CLTU_0_TC_Packet_Counter[2] , \CLTU_0_TC_Packet_Counter[3] , 
        \CLTU_0_TC_Packet_Counter[4] , \CLTU_0_TC_Packet_Counter[5] , 
        \CLTU_0_TC_Packet_Counter[6] , \CLTU_0_TC_Packet_Counter[7] , 
        \CLTU_0_TC_Packet_Counter[8] , \CLTU_0_TC_Packet_Counter[9] , 
        \CLTU_0_TC_Packet_Counter[10] , \CLTU_0_TC_Packet_Counter[11] , 
        \CLTU_0_TC_Packet_Counter[12] , \CLTU_0_TC_Packet_Counter[13] , 
        \CLTU_0_TC_Packet_Counter[14] , \CLTU_0_TC_Packet_Counter[15] , 
        \CLTU_0_TC_Packet_Counter[16] , \CLTU_0_TC_Packet_Counter[17] , 
        \CLTU_0_TC_Packet_Counter[18] , \CLTU_0_TC_Packet_Counter[19] , 
        \CLTU_0_TC_Packet_Counter[20] , \CLTU_0_TC_Packet_Counter[21] , 
        \CLTU_0_TC_Packet_Counter[22] , \CLTU_0_TC_Packet_Counter[23] , 
        \CLTU_0_TC_Packet_Counter[24] , \CLTU_0_TC_Packet_Counter[25] , 
        \CLTU_0_TC_Packet_Counter[26] , \CLTU_0_TC_Packet_Counter[27] , 
        \CLTU_0_TC_Packet_Counter[28] , \CLTU_0_TC_Packet_Counter[29] , 
        \CLTU_0_TC_Packet_Counter[30] , \CLTU_0_TC_Packet_Counter[31] , 
        \CLTU_0_TC_Error_Counter[1] , \CLTU_0_TC_Error_Counter[2] , 
        \CLTU_0_TC_Error_Counter[3] , \CLTU_0_TC_Error_Counter[4] , 
        \CLTU_0_TC_Error_Counter[5] , \CLTU_0_TC_Error_Counter[6] , 
        \CLTU_0_TC_Error_Counter[7] , \CLTU_0_TC_Error_Counter[8] , 
        \CLTU_0_TC_Error_Counter[9] , \CLTU_0_TC_Error_Counter[10] , 
        \CLTU_0_TC_Error_Counter[11] , \CLTU_0_TC_Error_Counter[12] , 
        \CLTU_0_TC_Error_Counter[13] , \CLTU_0_TC_Error_Counter[14] , 
        \CLTU_0_TC_Error_Counter[15] , \CLTU_0_TC_Error_Counter[16] , 
        \CLTU_0_TC_Error_Counter[17] , \CLTU_0_TC_Error_Counter[18] , 
        \CLTU_0_TC_Error_Counter[19] , \CLTU_0_TC_Error_Counter[20] , 
        \CLTU_0_TC_Error_Counter[21] , \CLTU_0_TC_Error_Counter[22] , 
        \CLTU_0_TC_Error_Counter[23] , \CLTU_0_TC_Error_Counter[24] , 
        \CLTU_0_TC_Error_Counter[25] , \CLTU_0_TC_Error_Counter[26] , 
        \CLTU_0_TC_Error_Counter[27] , \CLTU_0_TC_Error_Counter[28] , 
        \CLTU_0_TC_Error_Counter[29] , \CLTU_0_TC_Error_Counter[30] , 
        \CLTU_0_TC_Error_Counter[31] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[0] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[1] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[2] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[3] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[4] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[5] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[6] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[7] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[8] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[9] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[10] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[11] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[12] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[13] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[14] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[15] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[16] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[17] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[18] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[19] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[20] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[21] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[22] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[23] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[24] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[25] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[26] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[27] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[28] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[29] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[30] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[31] , 
        \divider_0.Bit_Count_16dec_i_1[3] , ENASM_i_0, N_623_i_0, 
        RX_GPIO1_ibuf_net_1, TX_GPIO1_ibuf_net_1;
    
    test_4463andcpuopration_MSS test_4463andcpuopration_MSS_0 (
        .CoreAPB3_0_APBmslave3_PADDR({
        \CoreAPB3_0_APBmslave3_PADDR[31] , 
        \CoreAPB3_0_APBmslave3_PADDR[30] , 
        \CoreAPB3_0_APBmslave3_PADDR[29] , 
        \CoreAPB3_0_APBmslave3_PADDR[28] , 
        \CoreAPB3_0_APBmslave3_PADDR[27] , 
        \CoreAPB3_0_APBmslave3_PADDR[26] , 
        \CoreAPB3_0_APBmslave3_PADDR[25] , 
        \CoreAPB3_0_APBmslave3_PADDR[24] , 
        \CoreAPB3_0_APBmslave3_PADDR[23] , 
        \CoreAPB3_0_APBmslave3_PADDR[22] , 
        \CoreAPB3_0_APBmslave3_PADDR[21] , 
        \CoreAPB3_0_APBmslave3_PADDR[20] , 
        \CoreAPB3_0_APBmslave3_PADDR[19] , 
        \CoreAPB3_0_APBmslave3_PADDR[18] , 
        \CoreAPB3_0_APBmslave3_PADDR[17] , 
        \CoreAPB3_0_APBmslave3_PADDR[16] , 
        \CoreAPB3_0_APBmslave3_PADDR[15] , 
        \CoreAPB3_0_APBmslave3_PADDR[14] , 
        \CoreAPB3_0_APBmslave3_PADDR[13] , 
        \CoreAPB3_0_APBmslave3_PADDR[12] , 
        \CoreAPB3_0_APBmslave3_PADDR[11] , 
        \CoreAPB3_0_APBmslave3_PADDR[10] , 
        \CoreAPB3_0_APBmslave3_PADDR[9] , 
        \CoreAPB3_0_APBmslave3_PADDR[8] , 
        \CoreAPB3_0_APBmslave3_PADDR[7] , 
        \CoreAPB3_0_APBmslave3_PADDR[6] , 
        \CoreAPB3_0_APBmslave3_PADDR[5] , 
        \CoreAPB3_0_APBmslave3_PADDR[4] , 
        \CoreAPB3_0_APBmslave3_PADDR[3] , 
        \CoreAPB3_0_APBmslave3_PADDR[2] , 
        \CoreAPB3_0_APBmslave3_PADDR[1] , 
        \CoreAPB3_0_APBmslave3_PADDR[0] }), 
        .CoreAPB3_0_APBmslave3_PWDATA({
        \CoreAPB3_0_APBmslave3_PWDATA[31] , 
        \CoreAPB3_0_APBmslave3_PWDATA[30] , 
        \CoreAPB3_0_APBmslave3_PWDATA[29] , 
        \CoreAPB3_0_APBmslave3_PWDATA[28] , 
        \CoreAPB3_0_APBmslave3_PWDATA[27] , 
        \CoreAPB3_0_APBmslave3_PWDATA[26] , 
        \CoreAPB3_0_APBmslave3_PWDATA[25] , 
        \CoreAPB3_0_APBmslave3_PWDATA[24] , 
        \CoreAPB3_0_APBmslave3_PWDATA[23] , 
        \CoreAPB3_0_APBmslave3_PWDATA[22] , 
        \CoreAPB3_0_APBmslave3_PWDATA[21] , 
        \CoreAPB3_0_APBmslave3_PWDATA[20] , 
        \CoreAPB3_0_APBmslave3_PWDATA[19] , 
        \CoreAPB3_0_APBmslave3_PWDATA[18] , 
        \CoreAPB3_0_APBmslave3_PWDATA[17] , 
        \CoreAPB3_0_APBmslave3_PWDATA[16] , 
        \CoreAPB3_0_APBmslave3_PWDATA[15] , 
        \CoreAPB3_0_APBmslave3_PWDATA[14] , 
        \CoreAPB3_0_APBmslave3_PWDATA[13] , 
        \CoreAPB3_0_APBmslave3_PWDATA[12] , 
        \CoreAPB3_0_APBmslave3_PWDATA[11] , 
        \CoreAPB3_0_APBmslave3_PWDATA[10] , 
        \CoreAPB3_0_APBmslave3_PWDATA[9] , 
        \CoreAPB3_0_APBmslave3_PWDATA[8] , 
        \CoreAPB3_0_APBmslave3_PWDATA[7] , 
        \CoreAPB3_0_APBmslave3_PWDATA[6] , 
        \CoreAPB3_0_APBmslave3_PWDATA[5] , 
        \CoreAPB3_0_APBmslave3_PWDATA[4] , 
        \CoreAPB3_0_APBmslave3_PWDATA[3] , 
        \CoreAPB3_0_APBmslave3_PWDATA[2] , 
        \CoreAPB3_0_APBmslave3_PWDATA[1] , 
        \CoreAPB3_0_APBmslave3_PWDATA[0] }), .Glue_Logic_0_Flag_Int_0({
        \Glue_Logic_0_Flag_Int_0[0] }), 
        .test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA({
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[31] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[30] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[29] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[28] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[27] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[26] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[25] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[24] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[23] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[22] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[21] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[20] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[19] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[18] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[17] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[16] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[0] }), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .SPI_CLK_c(
        SPI_CLK_c), .CAN1_RX_c(CAN1_RX_c), 
        .CoreAPB3_0_APBmslave3_PENABLE(CoreAPB3_0_APBmslave3_PENABLE), 
        .test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), 
        .CoreAPB3_0_APBmslave3_PWRITE(CoreAPB3_0_APBmslave3_PWRITE), 
        .SW_c(SW_c), .RX_SDN_c(RX_SDN_c), .Z3V_EN_c(\A3.3V_EN_c ), 
        .L4463_TX_CS_c(L4463_TX_CS_c), .L4463_RX_CS_c(L4463_RX_CS_c), 
        .TX_SDN_c(TX_SDN_c), .L3V3_EN1_c(L3V3_EN1_c), .ADC_CSTART_c(
        ADC_CSTART_c), .TXD4_c(TXD4_c), .SPI_FRAM_CS_c(SPI_FRAM_CS_c), 
        .SPI_MOSI_c(SPI_MOSI_c), .ADC_CS_c(ADC_CS_c), .ADC_FS_c(
        ADC_FS_c), .ADC_PWDN_c(ADC_PWDN_c), .L4V_EN_c(L4V_EN_c), 
        .ANT_SW1_c(ANT_SW1_c), 
        .test_4463andcpuopration_MSS_0_GPIO_15_M2F(
        test_4463andcpuopration_MSS_0_GPIO_15_M2F), .L3V3_EN2_c(
        L3V3_EN2_c), .CAN1_TX_c(CAN1_TX_c), .N_623_i_0(N_623_i_0), 
        .ADC_INT_c(ADC_INT_c), .L4V_PG_c(L4V_PG_c), .BOARD_NO_c(
        BOARD_NO_c), .RXD4_c(RXD4_c), .SPI_MISO_c(SPI_MISO_c), 
        .SYSRESET_0_POWER_ON_RESET_N(SYSRESET_0_POWER_ON_RESET_N), 
        .OSC_0_XTLOSC_O2F(OSC_0_XTLOSC_O2F));
    INBUF CCA_NIRQ_ibuf (.PAD(CCA_NIRQ), .Y(CCA_NIRQ_c));
    OUTBUF TX_SDN_obuf (.D(TX_SDN_c), .PAD(TX_SDN));
    Switch Switch_0 (.stream({\ASM_Generato_0.stream[0] }), .pn_reg({
        \Randomizer_0.pn_reg[0] }), .Switch_0_EnOut(Switch_0_EnOut), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .P_CLK(P_CLK), 
        .c_in(c_in), .ASM_OUT(ASM_OUT), .S_OUT_0(S_OUT_0), .P_OUT(
        P_OUT));
    CPU_W_HDL_R CPU_W_HDL_R_0 (.CPU_W_HDL_R_0_TM_Packet_Counter({
        \CPU_W_HDL_R_0_TM_Packet_Counter[31] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[30] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[29] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[28] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[27] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[26] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[25] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[24] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[23] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[22] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[21] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[20] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[19] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[18] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[17] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[16] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[15] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[14] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[13] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[12] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[11] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[10] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[9] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[8] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[7] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[6] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[5] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[4] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[3] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[2] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[1] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[0] }), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_9(\CPU_W_HDL_R_0_USER_RA_TRP1[9] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_0(\CPU_W_HDL_R_0_USER_RA_TRP1[0] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_1(\CPU_W_HDL_R_0_USER_RA_TRP1[1] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_2(\CPU_W_HDL_R_0_USER_RA_TRP1[2] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_3(\CPU_W_HDL_R_0_USER_RA_TRP1[3] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_4(\CPU_W_HDL_R_0_USER_RA_TRP1[4] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_5(\CPU_W_HDL_R_0_USER_RA_TRP1[5] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_6(\CPU_W_HDL_R_0_USER_RA_TRP1[6] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_7(\CPU_W_HDL_R_0_USER_RA_TRP1[7] ), 
        .ENASM(ENASM), .ENASM_i_0(ENASM_i_0), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .P_CLK(P_CLK), 
        .CPU_W_HDL_R_0_USER_REN_TRP1(CPU_W_HDL_R_0_USER_REN_TRP1), 
        .CPU_W_HDL_R_0_Flag_B_Tx_Finish(CPU_W_HDL_R_0_Flag_B_Tx_Finish)
        , .CPU_W_HDL_R_0_Flag_A_Tx_Finish(
        CPU_W_HDL_R_0_Flag_A_Tx_Finish), .ENCRC(ENCRC), 
        .Glue_Logic_0_Flag_B_Tx(Glue_Logic_0_Flag_B_Tx), .TXD4_net_0(
        TXD4_net_0), .pending(pending), .En_read_buff(En_read_buff));
    Randomizer Randomizer_0 (.pn_reg_0(\Randomizer_0.pn_reg[0] ), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .P_CLK(P_CLK), 
        .S_OUT_0(S_OUT_0));
    OUTBUF L3V3_EN1_obuf (.D(L3V3_EN1_c), .PAD(L3V3_EN1));
    OUTBUF L3V3_EN2_obuf (.D(L3V3_EN2_c), .PAD(L3V3_EN2));
    HDL_W_CPU_R_BUFF HDL_W_CPU_R_BUFF_0 (
        .HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1({
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[3] , 
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[2] , 
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[1] , 
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0] }), 
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1({
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[31] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[30] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[29] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[28] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[27] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[26] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[25] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[24] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[23] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[22] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[21] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[20] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[19] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[18] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[17] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[16] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[15] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[14] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[13] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[12] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[11] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[10] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[9] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[8] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[7] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[6] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[5] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[4] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[3] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[2] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[1] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[0] }), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .RX_GPIO1_c(
        RX_GPIO1_c), .EnIP(EnIP), 
        .HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish(
        HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish), 
        .HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish(
        HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish), 
        .HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1(
        HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1), .Glue_Logic_0_Flag_B_Rx(
        Glue_Logic_0_Flag_B_Rx), .Flag_RX(Flag_RX), .C_1(C_1), 
        .TC_Decode_0_IP_END_O(TC_Decode_0_IP_END_O), .FALG_FINISH_A_0(
        FALG_FINISH_A_0));
    DATA_OUT DATA_OUT_0 (.shift1_reg_4(
        \Convolutional_Encoder_0.shift1_reg[4] ), .shift1_reg_0(
        \Convolutional_Encoder_0.shift1_reg[0] ), .TX_GPIO0_c(
        TX_GPIO0_c), .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .TX_GPIO1_c(
        TX_GPIO1_c), .Convolutional_Encoder_out_1_0(
        \Convolutional_Encoder_0.Convolutional_Encoder_out_1_0 ), 
        .P_CLK(P_CLK));
    OUTBUF RX_SDN_obuf (.D(RX_SDN_c), .PAD(RX_SDN));
    OUTBUF CAN1_RX_obuf (.D(CAN1_RX_c), .PAD(CAN1_RX));
    INBUF RXD4_ibuf (.PAD(RXD4), .Y(RXD4_c));
    CoreAPB3_Z1 CoreAPB3_0 (.CoreAPB3_0_APBmslave3_PADDR({
        \CoreAPB3_0_APBmslave3_PADDR[31] , 
        \CoreAPB3_0_APBmslave3_PADDR[30] , 
        \CoreAPB3_0_APBmslave3_PADDR[29] , 
        \CoreAPB3_0_APBmslave3_PADDR[28] }), 
        .CoreAPB3_0_APBmslave3_PRDATA({
        \CoreAPB3_0_APBmslave3_PRDATA[31] , 
        \CoreAPB3_0_APBmslave3_PRDATA[30] , 
        \CoreAPB3_0_APBmslave3_PRDATA[29] , 
        \CoreAPB3_0_APBmslave3_PRDATA[28] , 
        \CoreAPB3_0_APBmslave3_PRDATA[27] , 
        \CoreAPB3_0_APBmslave3_PRDATA[26] , 
        \CoreAPB3_0_APBmslave3_PRDATA[25] , 
        \CoreAPB3_0_APBmslave3_PRDATA[24] , 
        \CoreAPB3_0_APBmslave3_PRDATA[23] , 
        \CoreAPB3_0_APBmslave3_PRDATA[22] , 
        \CoreAPB3_0_APBmslave3_PRDATA[21] , 
        \CoreAPB3_0_APBmslave3_PRDATA[20] , 
        \CoreAPB3_0_APBmslave3_PRDATA[19] , 
        \CoreAPB3_0_APBmslave3_PRDATA[18] , 
        \CoreAPB3_0_APBmslave3_PRDATA[17] , 
        \CoreAPB3_0_APBmslave3_PRDATA[16] , 
        \CoreAPB3_0_APBmslave3_PRDATA[15] , 
        \CoreAPB3_0_APBmslave3_PRDATA[14] , 
        \CoreAPB3_0_APBmslave3_PRDATA[13] , 
        \CoreAPB3_0_APBmslave3_PRDATA[12] , 
        \CoreAPB3_0_APBmslave3_PRDATA[11] , 
        \CoreAPB3_0_APBmslave3_PRDATA[10] , 
        \CoreAPB3_0_APBmslave3_PRDATA[9] , 
        \CoreAPB3_0_APBmslave3_PRDATA[8] , 
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] }), 
        .test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA({
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[31] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[30] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[29] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[28] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[27] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[26] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[25] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[24] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[23] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[22] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[21] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[20] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[19] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[18] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[17] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[16] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PRDATA[0] }), 
        .iPSELS_raw23(\CoreAPB3_0.iPSELS_raw23 ), 
        .test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), 
        .CoreAPB3_0_APBmslave3_PREADY(CoreAPB3_0_APBmslave3_PREADY), 
        .N_623_i_0(N_623_i_0));
    VCC VCC (.Y(VCC_net_1));
    test_4463andcpuopration_COREEDAC_1_COREEDAC_Z9 COREEDAC_1 (
        .HDL_W_CPU_R_BUFF_0_MSG_TRP1({
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[31] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[30] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[29] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[28] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[27] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[26] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[25] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[24] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[23] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[22] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[21] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[20] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[19] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[18] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[17] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[16] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[15] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[14] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[13] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[12] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[11] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[10] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[9] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[8] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[7] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[6] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[5] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[4] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[3] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[2] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[1] , 
        \HDL_W_CPU_R_BUFF_0_MSG_TRP1[0] }), .COREEDAC_1_DATA_OUT({
        \COREEDAC_1_DATA_OUT[31] , \COREEDAC_1_DATA_OUT[30] , 
        \COREEDAC_1_DATA_OUT[29] , \COREEDAC_1_DATA_OUT[28] , 
        \COREEDAC_1_DATA_OUT[27] , \COREEDAC_1_DATA_OUT[26] , 
        \COREEDAC_1_DATA_OUT[25] , \COREEDAC_1_DATA_OUT[24] , 
        \COREEDAC_1_DATA_OUT[23] , \COREEDAC_1_DATA_OUT[22] , 
        \COREEDAC_1_DATA_OUT[21] , \COREEDAC_1_DATA_OUT[20] , 
        \COREEDAC_1_DATA_OUT[19] , \COREEDAC_1_DATA_OUT[18] , 
        \COREEDAC_1_DATA_OUT[17] , \COREEDAC_1_DATA_OUT[16] , 
        \COREEDAC_1_DATA_OUT[15] , \COREEDAC_1_DATA_OUT[14] , 
        \COREEDAC_1_DATA_OUT[13] , \COREEDAC_1_DATA_OUT[12] , 
        \COREEDAC_1_DATA_OUT[11] , \COREEDAC_1_DATA_OUT[10] , 
        \COREEDAC_1_DATA_OUT[9] , \COREEDAC_1_DATA_OUT[8] , 
        \COREEDAC_1_DATA_OUT[7] , \COREEDAC_1_DATA_OUT[6] , 
        \COREEDAC_1_DATA_OUT[5] , \COREEDAC_1_DATA_OUT[4] , 
        \COREEDAC_1_DATA_OUT[3] , \COREEDAC_1_DATA_OUT[2] , 
        \COREEDAC_1_DATA_OUT[1] , \COREEDAC_1_DATA_OUT[0] }), 
        .Glue_Logic_0_USER_RA_TRP1_1({\Glue_Logic_0_USER_RA_TRP1_1[3] , 
        \Glue_Logic_0_USER_RA_TRP1_1[2] , 
        \Glue_Logic_0_USER_RA_TRP1_1[1] , 
        \Glue_Logic_0_USER_RA_TRP1_1[0] }), 
        .HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1({
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[3] , 
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[2] , 
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[1] , 
        \HDL_W_CPU_R_BUFF_0_MSG_WA_TRP1_1[0] }), .OSC_0_XTLOSC_O2F(
        OSC_0_XTLOSC_O2F), .Glue_Logic_0_USER_REN_TRP1(
        Glue_Logic_0_USER_REN_TRP1), .RX_GPIO1_c(RX_GPIO1_c), 
        .HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1(
        HDL_W_CPU_R_BUFF_0_USER_WEN_TRP1));
    divider divider_0 (.Bit_Count_16dec_i_1({
        \divider_0.Bit_Count_16dec_i_1[3] }), .P_CLK(P_CLK), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .TX_GPIO1_c(
        TX_GPIO1_c));
    INBUF BOARD_NO_ibuf (.PAD(BOARD_NO), .Y(BOARD_NO_c));
    OUTBUF SPI_FRAM_CS_obuf (.D(SPI_FRAM_CS_c), .PAD(SPI_FRAM_CS));
    OUTBUF ADC_CS_obuf (.D(ADC_CS_c), .PAD(ADC_CS));
    OUTBUF SPI_MOSI_obuf (.D(SPI_MOSI_c), .PAD(SPI_MOSI));
    INBUF SPI_MISO_ibuf (.PAD(SPI_MISO), .Y(SPI_MISO_c));
    test_4463andcpuopration_OSC_0_OSC OSC_0 (.OSC_0_XTLOSC_O2F(
        OSC_0_XTLOSC_O2F), .XTL(XTL));
    INBUF ADC_INT_ibuf (.PAD(ADC_INT), .Y(ADC_INT_c));
    OUTBUF ANT_SW1_obuf (.D(ANT_SW1_c), .PAD(ANT_SW1));
    INBUF RX_GPIO0_ibuf (.PAD(RX_GPIO0), .Y(RX_GPIO0_c));
    ASM_Generato ASM_Generato_0 (.stream_0(\ASM_Generato_0.stream[0] ), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .P_CLK(P_CLK), 
        .ASM_OUT(ASM_OUT), .pending(pending), .ENASM_i_0(ENASM_i_0), 
        .ENASM(ENASM));
    OR2 OR2_0 (.A(test_4463andcpuopration_MSS_0_GPIO_15_M2F), .B(
        GND_net_1), .Y(PA4V_ON_c));
    GND GND (.Y(GND_net_1));
    OUTBUF ADC_PWDN_obuf (.D(ADC_PWDN_c), .PAD(ADC_PWDN));
    OUTBUF ADC_FS_obuf (.D(ADC_FS_c), .PAD(ADC_FS));
    parallel_to_serial parallel_to_serial_0 (.TM_RSENC_0_CODEOUTP({
        \TM_RSENC_0_CODEOUTP[7] , \TM_RSENC_0_CODEOUTP[6] , 
        \TM_RSENC_0_CODEOUTP[5] , \TM_RSENC_0_CODEOUTP[4] , 
        \TM_RSENC_0_CODEOUTP[3] , \TM_RSENC_0_CODEOUTP[2] , 
        \TM_RSENC_0_CODEOUTP[1] , \TM_RSENC_0_CODEOUTP[0] }), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .P_CLK(P_CLK), 
        .S_OUT_0(S_OUT_0), .TM_RSENC_0_RDY(TM_RSENC_0_RDY), .P_OUT(
        P_OUT), .En_read_buff(En_read_buff));
    CLTU CLTU_0 (.CLTU_0_TC_Packet_Counter({
        \CLTU_0_TC_Packet_Counter[31] , \CLTU_0_TC_Packet_Counter[30] , 
        \CLTU_0_TC_Packet_Counter[29] , \CLTU_0_TC_Packet_Counter[28] , 
        \CLTU_0_TC_Packet_Counter[27] , \CLTU_0_TC_Packet_Counter[26] , 
        \CLTU_0_TC_Packet_Counter[25] , \CLTU_0_TC_Packet_Counter[24] , 
        \CLTU_0_TC_Packet_Counter[23] , \CLTU_0_TC_Packet_Counter[22] , 
        \CLTU_0_TC_Packet_Counter[21] , \CLTU_0_TC_Packet_Counter[20] , 
        \CLTU_0_TC_Packet_Counter[19] , \CLTU_0_TC_Packet_Counter[18] , 
        \CLTU_0_TC_Packet_Counter[17] , \CLTU_0_TC_Packet_Counter[16] , 
        \CLTU_0_TC_Packet_Counter[15] , \CLTU_0_TC_Packet_Counter[14] , 
        \CLTU_0_TC_Packet_Counter[13] , \CLTU_0_TC_Packet_Counter[12] , 
        \CLTU_0_TC_Packet_Counter[11] , \CLTU_0_TC_Packet_Counter[10] , 
        \CLTU_0_TC_Packet_Counter[9] , \CLTU_0_TC_Packet_Counter[8] , 
        \CLTU_0_TC_Packet_Counter[7] , \CLTU_0_TC_Packet_Counter[6] , 
        \CLTU_0_TC_Packet_Counter[5] , \CLTU_0_TC_Packet_Counter[4] , 
        \CLTU_0_TC_Packet_Counter[3] , \CLTU_0_TC_Packet_Counter[2] , 
        \CLTU_0_TC_Packet_Counter[1] , \CLTU_0_TC_Packet_Counter[0] }), 
        .CLTU_0_TC_Error_Counter({\CLTU_0_TC_Error_Counter[31] , 
        \CLTU_0_TC_Error_Counter[30] , \CLTU_0_TC_Error_Counter[29] , 
        \CLTU_0_TC_Error_Counter[28] , \CLTU_0_TC_Error_Counter[27] , 
        \CLTU_0_TC_Error_Counter[26] , \CLTU_0_TC_Error_Counter[25] , 
        \CLTU_0_TC_Error_Counter[24] , \CLTU_0_TC_Error_Counter[23] , 
        \CLTU_0_TC_Error_Counter[22] , \CLTU_0_TC_Error_Counter[21] , 
        \CLTU_0_TC_Error_Counter[20] , \CLTU_0_TC_Error_Counter[19] , 
        \CLTU_0_TC_Error_Counter[18] , \CLTU_0_TC_Error_Counter[17] , 
        \CLTU_0_TC_Error_Counter[16] , \CLTU_0_TC_Error_Counter[15] , 
        \CLTU_0_TC_Error_Counter[14] , \CLTU_0_TC_Error_Counter[13] , 
        \CLTU_0_TC_Error_Counter[12] , \CLTU_0_TC_Error_Counter[11] , 
        \CLTU_0_TC_Error_Counter[10] , \CLTU_0_TC_Error_Counter[9] , 
        \CLTU_0_TC_Error_Counter[8] , \CLTU_0_TC_Error_Counter[7] , 
        \CLTU_0_TC_Error_Counter[6] , \CLTU_0_TC_Error_Counter[5] , 
        \CLTU_0_TC_Error_Counter[4] , \CLTU_0_TC_Error_Counter[3] , 
        \CLTU_0_TC_Error_Counter[2] , \CLTU_0_TC_Error_Counter[1] , 
        \CLTU_0_TC_Error_Counter[0] }), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .RX_GPIO1_c(
        RX_GPIO1_c), .CLTU_0_IP_END(CLTU_0_IP_END), .A_1(A_1), 
        .ENASM_0(ENASM_0), .CLTU_0_Flag_RX_ing(CLTU_0_Flag_RX_ing), 
        .CLTU_0_Block_ErrO(CLTU_0_Block_ErrO), .CCA_NIRQ_c(CCA_NIRQ_c), 
        .RX_GPIO0_c(RX_GPIO0_c));
    OUTBUF CAN1_RS_obuf (.D(GND_net_1), .PAD(CAN1_RS));
    OUTBUF PA4V_ON_obuf (.D(PA4V_ON_c), .PAD(PA4V_ON));
    OUTBUF ANT_SW2_obuf (.D(ANT_SW2_c), .PAD(ANT_SW2));
    CLKINT RX_GPIO1_ibuf_RNIEM3F (.A(RX_GPIO1_ibuf_net_1), .Y(
        RX_GPIO1_c));
    CLKINT TX_GPIO1_ibuf_RNIGE8B (.A(TX_GPIO1_ibuf_net_1), .Y(
        TX_GPIO1_c));
    INBUF TX_GPIO1_ibuf (.PAD(TX_GPIO1), .Y(TX_GPIO1_ibuf_net_1));
    TM_RSENC TM_RSENC_0 (.Bit_Count_16dec_i_1({
        \divider_0.Bit_Count_16dec_i_1[3] }), .RSControl_0_DATAINP({
        \RSControl_0_DATAINP[7] , \RSControl_0_DATAINP[6] , 
        \RSControl_0_DATAINP[5] , \RSControl_0_DATAINP[4] , 
        \RSControl_0_DATAINP[3] , \RSControl_0_DATAINP[2] , 
        \RSControl_0_DATAINP[1] , \RSControl_0_DATAINP[0] }), 
        .TM_RSENC_0_CODEOUTP({\TM_RSENC_0_CODEOUTP[7] , 
        \TM_RSENC_0_CODEOUTP[6] , \TM_RSENC_0_CODEOUTP[5] , 
        \TM_RSENC_0_CODEOUTP[4] , \TM_RSENC_0_CODEOUTP[3] , 
        \TM_RSENC_0_CODEOUTP[2] , \TM_RSENC_0_CODEOUTP[1] , 
        \TM_RSENC_0_CODEOUTP[0] }), .TM_RSENC_0_RFD(TM_RSENC_0_RFD), 
        .RSControl_0_NGRST(RSControl_0_NGRST), .TM_RSENC_0_RFS(
        TM_RSENC_0_RFS), .RSControl_0_START(RSControl_0_START), 
        .TM_RSENC_0_RDY(TM_RSENC_0_RDY));
    OUTBUF SW_obuf (.D(SW_c), .PAD(SW));
    Glue_Logic_Z10 Glue_Logic_0 (.Glue_Logic_0_USER_RA_TRP1_1({
        \Glue_Logic_0_USER_RA_TRP1_1[3] , 
        \Glue_Logic_0_USER_RA_TRP1_1[2] , 
        \Glue_Logic_0_USER_RA_TRP1_1[1] , 
        \Glue_Logic_0_USER_RA_TRP1_1[0] }), .Glue_Logic_0_MSG_WA_TRP1({
        \Glue_Logic_0_MSG_WA_TRP1[9] , \Glue_Logic_0_MSG_WA_TRP1[8] , 
        \Glue_Logic_0_MSG_WA_TRP1[7] , \Glue_Logic_0_MSG_WA_TRP1[6] , 
        \Glue_Logic_0_MSG_WA_TRP1[5] , \Glue_Logic_0_MSG_WA_TRP1[4] , 
        \Glue_Logic_0_MSG_WA_TRP1[3] , \Glue_Logic_0_MSG_WA_TRP1[2] , 
        \Glue_Logic_0_MSG_WA_TRP1[1] , \Glue_Logic_0_MSG_WA_TRP1[0] }), 
        .CoreAPB3_0_APBmslave3_PRDATA({
        \CoreAPB3_0_APBmslave3_PRDATA[31] , 
        \CoreAPB3_0_APBmslave3_PRDATA[30] , 
        \CoreAPB3_0_APBmslave3_PRDATA[29] , 
        \CoreAPB3_0_APBmslave3_PRDATA[28] , 
        \CoreAPB3_0_APBmslave3_PRDATA[27] , 
        \CoreAPB3_0_APBmslave3_PRDATA[26] , 
        \CoreAPB3_0_APBmslave3_PRDATA[25] , 
        \CoreAPB3_0_APBmslave3_PRDATA[24] , 
        \CoreAPB3_0_APBmslave3_PRDATA[23] , 
        \CoreAPB3_0_APBmslave3_PRDATA[22] , 
        \CoreAPB3_0_APBmslave3_PRDATA[21] , 
        \CoreAPB3_0_APBmslave3_PRDATA[20] , 
        \CoreAPB3_0_APBmslave3_PRDATA[19] , 
        \CoreAPB3_0_APBmslave3_PRDATA[18] , 
        \CoreAPB3_0_APBmslave3_PRDATA[17] , 
        \CoreAPB3_0_APBmslave3_PRDATA[16] , 
        \CoreAPB3_0_APBmslave3_PRDATA[15] , 
        \CoreAPB3_0_APBmslave3_PRDATA[14] , 
        \CoreAPB3_0_APBmslave3_PRDATA[13] , 
        \CoreAPB3_0_APBmslave3_PRDATA[12] , 
        \CoreAPB3_0_APBmslave3_PRDATA[11] , 
        \CoreAPB3_0_APBmslave3_PRDATA[10] , 
        \CoreAPB3_0_APBmslave3_PRDATA[9] , 
        \CoreAPB3_0_APBmslave3_PRDATA[8] , 
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] }), .Glue_Logic_0_MSG_TRP1({
        \Glue_Logic_0_MSG_TRP1[7] , \Glue_Logic_0_MSG_TRP1[6] , 
        \Glue_Logic_0_MSG_TRP1[5] , \Glue_Logic_0_MSG_TRP1[4] , 
        \Glue_Logic_0_MSG_TRP1[3] , \Glue_Logic_0_MSG_TRP1[2] , 
        \Glue_Logic_0_MSG_TRP1[1] , \Glue_Logic_0_MSG_TRP1[0] }), 
        .Glue_Logic_0_Flag_Int_0({\Glue_Logic_0_Flag_Int_0[0] }), 
        .CoreAPB3_0_APBmslave3_PADDR({
        \CoreAPB3_0_APBmslave3_PADDR[31] , 
        \CoreAPB3_0_APBmslave3_PADDR[30] , 
        \CoreAPB3_0_APBmslave3_PADDR[29] , 
        \CoreAPB3_0_APBmslave3_PADDR[28] , 
        \CoreAPB3_0_APBmslave3_PADDR[27] , 
        \CoreAPB3_0_APBmslave3_PADDR[26] , 
        \CoreAPB3_0_APBmslave3_PADDR[25] , 
        \CoreAPB3_0_APBmslave3_PADDR[24] , 
        \CoreAPB3_0_APBmslave3_PADDR[23] , 
        \CoreAPB3_0_APBmslave3_PADDR[22] , 
        \CoreAPB3_0_APBmslave3_PADDR[21] , 
        \CoreAPB3_0_APBmslave3_PADDR[20] , 
        \CoreAPB3_0_APBmslave3_PADDR[19] , 
        \CoreAPB3_0_APBmslave3_PADDR[18] , 
        \CoreAPB3_0_APBmslave3_PADDR[17] , 
        \CoreAPB3_0_APBmslave3_PADDR[16] , 
        \CoreAPB3_0_APBmslave3_PADDR[15] , 
        \CoreAPB3_0_APBmslave3_PADDR[14] , 
        \CoreAPB3_0_APBmslave3_PADDR[13] , 
        \CoreAPB3_0_APBmslave3_PADDR[12] , 
        \CoreAPB3_0_APBmslave3_PADDR[11] , 
        \CoreAPB3_0_APBmslave3_PADDR[10] , 
        \CoreAPB3_0_APBmslave3_PADDR[9] , 
        \CoreAPB3_0_APBmslave3_PADDR[8] , 
        \CoreAPB3_0_APBmslave3_PADDR[7] , 
        \CoreAPB3_0_APBmslave3_PADDR[6] , 
        \CoreAPB3_0_APBmslave3_PADDR[5] , 
        \CoreAPB3_0_APBmslave3_PADDR[4] , 
        \CoreAPB3_0_APBmslave3_PADDR[3] , 
        \CoreAPB3_0_APBmslave3_PADDR[2] , 
        \CoreAPB3_0_APBmslave3_PADDR[1] , 
        \CoreAPB3_0_APBmslave3_PADDR[0] }), 
        .CoreAPB3_0_APBmslave3_PWDATA({
        \CoreAPB3_0_APBmslave3_PWDATA[31] , 
        \CoreAPB3_0_APBmslave3_PWDATA[30] , 
        \CoreAPB3_0_APBmslave3_PWDATA[29] , 
        \CoreAPB3_0_APBmslave3_PWDATA[28] , 
        \CoreAPB3_0_APBmslave3_PWDATA[27] , 
        \CoreAPB3_0_APBmslave3_PWDATA[26] , 
        \CoreAPB3_0_APBmslave3_PWDATA[25] , 
        \CoreAPB3_0_APBmslave3_PWDATA[24] , 
        \CoreAPB3_0_APBmslave3_PWDATA[23] , 
        \CoreAPB3_0_APBmslave3_PWDATA[22] , 
        \CoreAPB3_0_APBmslave3_PWDATA[21] , 
        \CoreAPB3_0_APBmslave3_PWDATA[20] , 
        \CoreAPB3_0_APBmslave3_PWDATA[19] , 
        \CoreAPB3_0_APBmslave3_PWDATA[18] , 
        \CoreAPB3_0_APBmslave3_PWDATA[17] , 
        \CoreAPB3_0_APBmslave3_PWDATA[16] , 
        \CoreAPB3_0_APBmslave3_PWDATA[15] , 
        \CoreAPB3_0_APBmslave3_PWDATA[14] , 
        \CoreAPB3_0_APBmslave3_PWDATA[13] , 
        \CoreAPB3_0_APBmslave3_PWDATA[12] , 
        \CoreAPB3_0_APBmslave3_PWDATA[11] , 
        \CoreAPB3_0_APBmslave3_PWDATA[10] , 
        \CoreAPB3_0_APBmslave3_PWDATA[9] , 
        \CoreAPB3_0_APBmslave3_PWDATA[8] , 
        \CoreAPB3_0_APBmslave3_PWDATA[7] , 
        \CoreAPB3_0_APBmslave3_PWDATA[6] , 
        \CoreAPB3_0_APBmslave3_PWDATA[5] , 
        \CoreAPB3_0_APBmslave3_PWDATA[4] , 
        \CoreAPB3_0_APBmslave3_PWDATA[3] , 
        \CoreAPB3_0_APBmslave3_PWDATA[2] , 
        \CoreAPB3_0_APBmslave3_PWDATA[1] , 
        \CoreAPB3_0_APBmslave3_PWDATA[0] }), 
        .CPU_W_HDL_R_0_TM_Packet_Counter({
        \CPU_W_HDL_R_0_TM_Packet_Counter[31] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[30] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[29] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[28] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[27] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[26] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[25] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[24] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[23] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[22] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[21] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[20] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[19] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[18] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[17] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[16] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[15] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[14] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[13] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[12] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[11] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[10] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[9] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[8] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[7] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[6] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[5] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[4] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[3] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[2] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[1] , 
        \CPU_W_HDL_R_0_TM_Packet_Counter[0] }), 
        .CLTU_0_TC_Packet_Counter({\CLTU_0_TC_Packet_Counter[31] , 
        \CLTU_0_TC_Packet_Counter[30] , \CLTU_0_TC_Packet_Counter[29] , 
        \CLTU_0_TC_Packet_Counter[28] , \CLTU_0_TC_Packet_Counter[27] , 
        \CLTU_0_TC_Packet_Counter[26] , \CLTU_0_TC_Packet_Counter[25] , 
        \CLTU_0_TC_Packet_Counter[24] , \CLTU_0_TC_Packet_Counter[23] , 
        \CLTU_0_TC_Packet_Counter[22] , \CLTU_0_TC_Packet_Counter[21] , 
        \CLTU_0_TC_Packet_Counter[20] , \CLTU_0_TC_Packet_Counter[19] , 
        \CLTU_0_TC_Packet_Counter[18] , \CLTU_0_TC_Packet_Counter[17] , 
        \CLTU_0_TC_Packet_Counter[16] , \CLTU_0_TC_Packet_Counter[15] , 
        \CLTU_0_TC_Packet_Counter[14] , \CLTU_0_TC_Packet_Counter[13] , 
        \CLTU_0_TC_Packet_Counter[12] , \CLTU_0_TC_Packet_Counter[11] , 
        \CLTU_0_TC_Packet_Counter[10] , \CLTU_0_TC_Packet_Counter[9] , 
        \CLTU_0_TC_Packet_Counter[8] , \CLTU_0_TC_Packet_Counter[7] , 
        \CLTU_0_TC_Packet_Counter[6] , \CLTU_0_TC_Packet_Counter[5] , 
        \CLTU_0_TC_Packet_Counter[4] , \CLTU_0_TC_Packet_Counter[3] , 
        \CLTU_0_TC_Packet_Counter[2] , \CLTU_0_TC_Packet_Counter[1] , 
        \CLTU_0_TC_Packet_Counter[0] }), .CLTU_0_TC_Error_Counter({
        \CLTU_0_TC_Error_Counter[31] , \CLTU_0_TC_Error_Counter[30] , 
        \CLTU_0_TC_Error_Counter[29] , \CLTU_0_TC_Error_Counter[28] , 
        \CLTU_0_TC_Error_Counter[27] , \CLTU_0_TC_Error_Counter[26] , 
        \CLTU_0_TC_Error_Counter[25] , \CLTU_0_TC_Error_Counter[24] , 
        \CLTU_0_TC_Error_Counter[23] , \CLTU_0_TC_Error_Counter[22] , 
        \CLTU_0_TC_Error_Counter[21] , \CLTU_0_TC_Error_Counter[20] , 
        \CLTU_0_TC_Error_Counter[19] , \CLTU_0_TC_Error_Counter[18] , 
        \CLTU_0_TC_Error_Counter[17] , \CLTU_0_TC_Error_Counter[16] , 
        \CLTU_0_TC_Error_Counter[15] , \CLTU_0_TC_Error_Counter[14] , 
        \CLTU_0_TC_Error_Counter[13] , \CLTU_0_TC_Error_Counter[12] , 
        \CLTU_0_TC_Error_Counter[11] , \CLTU_0_TC_Error_Counter[10] , 
        \CLTU_0_TC_Error_Counter[9] , \CLTU_0_TC_Error_Counter[8] , 
        \CLTU_0_TC_Error_Counter[7] , \CLTU_0_TC_Error_Counter[6] , 
        \CLTU_0_TC_Error_Counter[5] , \CLTU_0_TC_Error_Counter[4] , 
        \CLTU_0_TC_Error_Counter[3] , \CLTU_0_TC_Error_Counter[2] , 
        \CLTU_0_TC_Error_Counter[1] , \CLTU_0_TC_Error_Counter[0] }), 
        .COREEDAC_1_DATA_OUT({\COREEDAC_1_DATA_OUT[31] , 
        \COREEDAC_1_DATA_OUT[30] , \COREEDAC_1_DATA_OUT[29] , 
        \COREEDAC_1_DATA_OUT[28] , \COREEDAC_1_DATA_OUT[27] , 
        \COREEDAC_1_DATA_OUT[26] , \COREEDAC_1_DATA_OUT[25] , 
        \COREEDAC_1_DATA_OUT[24] , \COREEDAC_1_DATA_OUT[23] , 
        \COREEDAC_1_DATA_OUT[22] , \COREEDAC_1_DATA_OUT[21] , 
        \COREEDAC_1_DATA_OUT[20] , \COREEDAC_1_DATA_OUT[19] , 
        \COREEDAC_1_DATA_OUT[18] , \COREEDAC_1_DATA_OUT[17] , 
        \COREEDAC_1_DATA_OUT[16] , \COREEDAC_1_DATA_OUT[15] , 
        \COREEDAC_1_DATA_OUT[14] , \COREEDAC_1_DATA_OUT[13] , 
        \COREEDAC_1_DATA_OUT[12] , \COREEDAC_1_DATA_OUT[11] , 
        \COREEDAC_1_DATA_OUT[10] , \COREEDAC_1_DATA_OUT[9] , 
        \COREEDAC_1_DATA_OUT[8] , \COREEDAC_1_DATA_OUT[7] , 
        \COREEDAC_1_DATA_OUT[6] , \COREEDAC_1_DATA_OUT[5] , 
        \COREEDAC_1_DATA_OUT[4] , \COREEDAC_1_DATA_OUT[3] , 
        \COREEDAC_1_DATA_OUT[2] , \COREEDAC_1_DATA_OUT[1] , 
        \COREEDAC_1_DATA_OUT[0] }), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .OSC_0_XTLOSC_O2F(
        OSC_0_XTLOSC_O2F), .Glue_Logic_0_USER_REN_TRP1(
        Glue_Logic_0_USER_REN_TRP1), .Glue_Logic_0_Flag_B_Tx(
        Glue_Logic_0_Flag_B_Tx), .Glue_Logic_0_Flag_B_Rx(
        Glue_Logic_0_Flag_B_Rx), .TXD4_net_0(TXD4_net_0), .Flag_RX(
        Flag_RX), .Glue_Logic_0_USER_WEN_TRP1(
        Glue_Logic_0_USER_WEN_TRP1), .CoreAPB3_0_APBmslave3_PREADY(
        CoreAPB3_0_APBmslave3_PREADY), 
        .HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish(
        HDL_W_CPU_R_BUFF_0_Flag_A_HDL_Rec_Finish), 
        .CPU_W_HDL_R_0_Flag_A_Tx_Finish(CPU_W_HDL_R_0_Flag_A_Tx_Finish)
        , .HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish(
        HDL_W_CPU_R_BUFF_0_Flag_B_HDL_Rec_Finish), 
        .CPU_W_HDL_R_0_Flag_B_Tx_Finish(CPU_W_HDL_R_0_Flag_B_Tx_Finish)
        , .CoreAPB3_0_APBmslave3_PWRITE(CoreAPB3_0_APBmslave3_PWRITE), 
        .Switch_0_EnOut(Switch_0_EnOut), .CLTU_0_Flag_RX_ing(
        CLTU_0_Flag_RX_ing), 
        .test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx(
        test_4463andcpuopration_MSS_0_FIC_0_APB_MASTER_PSELx), 
        .CoreAPB3_0_APBmslave3_PENABLE(CoreAPB3_0_APBmslave3_PENABLE), 
        .iPSELS_raw23(\CoreAPB3_0.iPSELS_raw23 ));
    OUTBUF ADC_CSTART_obuf (.D(ADC_CSTART_c), .PAD(ADC_CSTART));
    OUTBUF \A3.3V_EN_obuf  (.D(\A3.3V_EN_c ), .PAD(\A3.3V_EN ));
    INBUF L4V_PG_ibuf (.PAD(L4V_PG), .Y(L4V_PG_c));
    OUTBUF L4463_TX_CS_obuf (.D(L4463_TX_CS_c), .PAD(L4463_TX_CS));
    OUTBUF SPI_CLK_obuf (.D(SPI_CLK_c), .PAD(SPI_CLK));
    OUTBUF L4V_EN_obuf (.D(L4V_EN_c), .PAD(L4V_EN));
    OUTBUF L4463_RX_CS_obuf (.D(L4463_RX_CS_c), .PAD(L4463_RX_CS));
    OUTBUF TX_GPIO0_obuf (.D(TX_GPIO0_c), .PAD(TX_GPIO0));
    INBUF RX_GPIO1_ibuf (.PAD(RX_GPIO1), .Y(RX_GPIO1_ibuf_net_1));
    OUTBUF TXD4_obuf (.D(TXD4_c), .PAD(TXD4));
    INV INV_0 (.A(ANT_SW1_c), .Y(ANT_SW2_c));
    Convolutional_Encoder Convolutional_Encoder_0 (.shift1_reg_4(
        \Convolutional_Encoder_0.shift1_reg[4] ), .shift1_reg_0(
        \Convolutional_Encoder_0.shift1_reg[0] ), 
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .P_CLK(P_CLK), 
        .c_in(c_in), .Convolutional_Encoder_out_1_0(
        \Convolutional_Encoder_0.Convolutional_Encoder_out_1_0 ));
    test_4463andcpuopration_COREEDAC_0_COREEDAC_Z5 COREEDAC_0 (
        .Glue_Logic_0_MSG_TRP1({\Glue_Logic_0_MSG_TRP1[7] , 
        \Glue_Logic_0_MSG_TRP1[6] , \Glue_Logic_0_MSG_TRP1[5] , 
        \Glue_Logic_0_MSG_TRP1[4] , \Glue_Logic_0_MSG_TRP1[3] , 
        \Glue_Logic_0_MSG_TRP1[2] , \Glue_Logic_0_MSG_TRP1[1] , 
        \Glue_Logic_0_MSG_TRP1[0] }), .CPU_W_HDL_R_0_DataO({
        \CPU_W_HDL_R_0_DataO[7] , \CPU_W_HDL_R_0_DataO[6] , 
        \CPU_W_HDL_R_0_DataO[5] , \CPU_W_HDL_R_0_DataO[4] , 
        \CPU_W_HDL_R_0_DataO[3] , \CPU_W_HDL_R_0_DataO[2] , 
        \CPU_W_HDL_R_0_DataO[1] , \CPU_W_HDL_R_0_DataO[0] }), 
        .Bit_Count_16dec_i_1({\divider_0.Bit_Count_16dec_i_1[3] }), 
        .Glue_Logic_0_MSG_WA_TRP1({\Glue_Logic_0_MSG_WA_TRP1[9] , 
        \Glue_Logic_0_MSG_WA_TRP1[8] , \Glue_Logic_0_MSG_WA_TRP1[7] , 
        \Glue_Logic_0_MSG_WA_TRP1[6] , \Glue_Logic_0_MSG_WA_TRP1[5] , 
        \Glue_Logic_0_MSG_WA_TRP1[4] , \Glue_Logic_0_MSG_WA_TRP1[3] , 
        \Glue_Logic_0_MSG_WA_TRP1[2] , \Glue_Logic_0_MSG_WA_TRP1[1] , 
        \Glue_Logic_0_MSG_WA_TRP1[0] }), .CPU_W_HDL_R_0_USER_RA_TRP1_0(
        \CPU_W_HDL_R_0_USER_RA_TRP1[0] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_1(\CPU_W_HDL_R_0_USER_RA_TRP1[1] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_2(\CPU_W_HDL_R_0_USER_RA_TRP1[2] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_3(\CPU_W_HDL_R_0_USER_RA_TRP1[3] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_4(\CPU_W_HDL_R_0_USER_RA_TRP1[4] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_5(\CPU_W_HDL_R_0_USER_RA_TRP1[5] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_6(\CPU_W_HDL_R_0_USER_RA_TRP1[6] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_7(\CPU_W_HDL_R_0_USER_RA_TRP1[7] ), 
        .CPU_W_HDL_R_0_USER_RA_TRP1_9(\CPU_W_HDL_R_0_USER_RA_TRP1[9] ), 
        .CPU_W_HDL_R_0_USER_REN_TRP1(CPU_W_HDL_R_0_USER_REN_TRP1), 
        .OSC_0_XTLOSC_O2F(OSC_0_XTLOSC_O2F), 
        .Glue_Logic_0_USER_WEN_TRP1(Glue_Logic_0_USER_WEN_TRP1));
    RSControl RSControl_0 (.Bit_Count_16dec_i_1({
        \divider_0.Bit_Count_16dec_i_1[3] }), .RSControl_0_DATAINP({
        \RSControl_0_DATAINP[7] , \RSControl_0_DATAINP[6] , 
        \RSControl_0_DATAINP[5] , \RSControl_0_DATAINP[4] , 
        \RSControl_0_DATAINP[3] , \RSControl_0_DATAINP[2] , 
        \RSControl_0_DATAINP[1] , \RSControl_0_DATAINP[0] }), 
        .CPU_W_HDL_R_0_DataO({\CPU_W_HDL_R_0_DataO[7] , 
        \CPU_W_HDL_R_0_DataO[6] , \CPU_W_HDL_R_0_DataO[5] , 
        \CPU_W_HDL_R_0_DataO[4] , \CPU_W_HDL_R_0_DataO[3] , 
        \CPU_W_HDL_R_0_DataO[2] , \CPU_W_HDL_R_0_DataO[1] , 
        \CPU_W_HDL_R_0_DataO[0] }), .RSControl_0_NGRST(
        RSControl_0_NGRST), .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .RSControl_0_START(
        RSControl_0_START), .TM_RSENC_0_RFD(TM_RSENC_0_RFD), .ENCRC(
        ENCRC), .TM_RSENC_0_RFS(TM_RSENC_0_RFS));
    SYSRESET SYSRESET_0 (.POWER_ON_RESET_N(SYSRESET_0_POWER_ON_RESET_N)
        , .DEVRST_N(DEVRST_N));
    INBUF CAN1_TX_ibuf (.PAD(CAN1_TX), .Y(CAN1_TX_c));
    TC_Decode TC_Decode_0 (.test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .RX_GPIO1_c(
        RX_GPIO1_c), .C_1(C_1), .FALG_FINISH_A_0(FALG_FINISH_A_0), 
        .TC_Decode_0_IP_END_O(TC_Decode_0_IP_END_O), .EnIP(EnIP), 
        .RXRandomize_0_Block_ErrO(RXRandomize_0_Block_ErrO), 
        .pending_0(pending_0), .ENCRC_0(ENCRC_0), 
        .RXRandomize_0_IP_END_O(RXRandomize_0_IP_END_O));
    OUTBUF CAN2_RS_obuf (.D(VCC_net_1), .PAD(CAN2_RS));
    RXRandomize RXRandomize_0 (
        .test_4463andcpuopration_MSS_0_GPIO_1_M2F(
        test_4463andcpuopration_MSS_0_GPIO_1_M2F), .RX_GPIO1_c(
        RX_GPIO1_c), .ENCRC_0(ENCRC_0), .pending_0(pending_0), 
        .RXRandomize_0_Block_ErrO(RXRandomize_0_Block_ErrO), 
        .CLTU_0_Block_ErrO(CLTU_0_Block_ErrO), .RXRandomize_0_IP_END_O(
        RXRandomize_0_IP_END_O), .CLTU_0_IP_END(CLTU_0_IP_END), 
        .ENASM_0(ENASM_0), .A_1(A_1));
    
endmodule
