// Copyright 2008 Actel Corporation. All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// 
// Revision: 0.2 April 30, 2008

// This is an automatically generated file

 `timescale 1 ns/100 ps

// Shortened Hamming code (13, 8) table-based encoder
// Use to generate non-synthesizable golden code 

  module bhv_enc_vlog (msg, coded); 
      input [7:0] msg; 
      output reg[12:0] coded; 
    always @ (msg) 
      case (msg) 
             0 : coded = 13'b0000000000000;   // 0 
             1 : coded = 13'b0000000100111;   // 39 
             2 : coded = 13'b0000001011001;   // 89 
             3 : coded = 13'b0000001111110;   // 126 
             4 : coded = 13'b0000010001110;   // 142 
             5 : coded = 13'b0000010101001;   // 169 
             6 : coded = 13'b0000011010111;   // 215 
             7 : coded = 13'b0000011110000;   // 240 
             8 : coded = 13'b0000100010011;   // 275 
             9 : coded = 13'b0000100110100;   // 308 
            10 : coded = 13'b0000101001010;   // 330 
            11 : coded = 13'b0000101101101;   // 365 
            12 : coded = 13'b0000110011101;   // 413 
            13 : coded = 13'b0000110111010;   // 442 
            14 : coded = 13'b0000111000100;   // 452 
            15 : coded = 13'b0000111100011;   // 483 
            16 : coded = 13'b0001000011100;   // 540 
            17 : coded = 13'b0001000111011;   // 571 
            18 : coded = 13'b0001001000101;   // 581 
            19 : coded = 13'b0001001100010;   // 610 
            20 : coded = 13'b0001010010010;   // 658 
            21 : coded = 13'b0001010110101;   // 693 
            22 : coded = 13'b0001011001011;   // 715 
            23 : coded = 13'b0001011101100;   // 748 
            24 : coded = 13'b0001100001111;   // 783 
            25 : coded = 13'b0001100101000;   // 808 
            26 : coded = 13'b0001101010110;   // 854 
            27 : coded = 13'b0001101110001;   // 881 
            28 : coded = 13'b0001110000001;   // 897 
            29 : coded = 13'b0001110100110;   // 934 
            30 : coded = 13'b0001111011000;   // 984 
            31 : coded = 13'b0001111111111;   // 1023 
            32 : coded = 13'b0010000001011;   // 1035 
            33 : coded = 13'b0010000101100;   // 1068 
            34 : coded = 13'b0010001010010;   // 1106 
            35 : coded = 13'b0010001110101;   // 1141 
            36 : coded = 13'b0010010000101;   // 1157 
            37 : coded = 13'b0010010100010;   // 1186 
            38 : coded = 13'b0010011011100;   // 1244 
            39 : coded = 13'b0010011111011;   // 1275 
            40 : coded = 13'b0010100011000;   // 1304 
            41 : coded = 13'b0010100111111;   // 1343 
            42 : coded = 13'b0010101000001;   // 1345 
            43 : coded = 13'b0010101100110;   // 1382 
            44 : coded = 13'b0010110010110;   // 1430 
            45 : coded = 13'b0010110110001;   // 1457 
            46 : coded = 13'b0010111001111;   // 1487 
            47 : coded = 13'b0010111101000;   // 1512 
            48 : coded = 13'b0011000010111;   // 1559 
            49 : coded = 13'b0011000110000;   // 1584 
            50 : coded = 13'b0011001001110;   // 1614 
            51 : coded = 13'b0011001101001;   // 1641 
            52 : coded = 13'b0011010011001;   // 1689 
            53 : coded = 13'b0011010111110;   // 1726 
            54 : coded = 13'b0011011000000;   // 1728 
            55 : coded = 13'b0011011100111;   // 1767 
            56 : coded = 13'b0011100000100;   // 1796 
            57 : coded = 13'b0011100100011;   // 1827 
            58 : coded = 13'b0011101011101;   // 1885 
            59 : coded = 13'b0011101111010;   // 1914 
            60 : coded = 13'b0011110001010;   // 1930 
            61 : coded = 13'b0011110101101;   // 1965 
            62 : coded = 13'b0011111010011;   // 2003 
            63 : coded = 13'b0011111110100;   // 2036 
            64 : coded = 13'b0100000010101;   // 2069 
            65 : coded = 13'b0100000110010;   // 2098 
            66 : coded = 13'b0100001001100;   // 2124 
            67 : coded = 13'b0100001101011;   // 2155 
            68 : coded = 13'b0100010011011;   // 2203 
            69 : coded = 13'b0100010111100;   // 2236 
            70 : coded = 13'b0100011000010;   // 2242 
            71 : coded = 13'b0100011100101;   // 2277 
            72 : coded = 13'b0100100000110;   // 2310 
            73 : coded = 13'b0100100100001;   // 2337 
            74 : coded = 13'b0100101011111;   // 2399 
            75 : coded = 13'b0100101111000;   // 2424 
            76 : coded = 13'b0100110001000;   // 2440 
            77 : coded = 13'b0100110101111;   // 2479 
            78 : coded = 13'b0100111010001;   // 2513 
            79 : coded = 13'b0100111110110;   // 2550 
            80 : coded = 13'b0101000001001;   // 2569 
            81 : coded = 13'b0101000101110;   // 2606 
            82 : coded = 13'b0101001010000;   // 2640 
            83 : coded = 13'b0101001110111;   // 2679 
            84 : coded = 13'b0101010000111;   // 2695 
            85 : coded = 13'b0101010100000;   // 2720 
            86 : coded = 13'b0101011011110;   // 2782 
            87 : coded = 13'b0101011111001;   // 2809 
            88 : coded = 13'b0101100011010;   // 2842 
            89 : coded = 13'b0101100111101;   // 2877 
            90 : coded = 13'b0101101000011;   // 2883 
            91 : coded = 13'b0101101100100;   // 2916 
            92 : coded = 13'b0101110010100;   // 2964 
            93 : coded = 13'b0101110110011;   // 2995 
            94 : coded = 13'b0101111001101;   // 3021 
            95 : coded = 13'b0101111101010;   // 3050 
            96 : coded = 13'b0110000011110;   // 3102 
            97 : coded = 13'b0110000111001;   // 3129 
            98 : coded = 13'b0110001000111;   // 3143 
            99 : coded = 13'b0110001100000;   // 3168 
           100 : coded = 13'b0110010010000;   // 3216 
           101 : coded = 13'b0110010110111;   // 3255 
           102 : coded = 13'b0110011001001;   // 3273 
           103 : coded = 13'b0110011101110;   // 3310 
           104 : coded = 13'b0110100001101;   // 3341 
           105 : coded = 13'b0110100101010;   // 3370 
           106 : coded = 13'b0110101010100;   // 3412 
           107 : coded = 13'b0110101110011;   // 3443 
           108 : coded = 13'b0110110000011;   // 3459 
           109 : coded = 13'b0110110100100;   // 3492 
           110 : coded = 13'b0110111011010;   // 3546 
           111 : coded = 13'b0110111111101;   // 3581 
           112 : coded = 13'b0111000000010;   // 3586 
           113 : coded = 13'b0111000100101;   // 3621 
           114 : coded = 13'b0111001011011;   // 3675 
           115 : coded = 13'b0111001111100;   // 3708 
           116 : coded = 13'b0111010001100;   // 3724 
           117 : coded = 13'b0111010101011;   // 3755 
           118 : coded = 13'b0111011010101;   // 3797 
           119 : coded = 13'b0111011110010;   // 3826 
           120 : coded = 13'b0111100010001;   // 3857 
           121 : coded = 13'b0111100110110;   // 3894 
           122 : coded = 13'b0111101001000;   // 3912 
           123 : coded = 13'b0111101101111;   // 3951 
           124 : coded = 13'b0111110011111;   // 3999 
           125 : coded = 13'b0111110111000;   // 4024 
           126 : coded = 13'b0111111000110;   // 4038 
           127 : coded = 13'b0111111100001;   // 4065 
           128 : coded = 13'b1000000010110;   // 4118 
           129 : coded = 13'b1000000110001;   // 4145 
           130 : coded = 13'b1000001001111;   // 4175 
           131 : coded = 13'b1000001101000;   // 4200 
           132 : coded = 13'b1000010011000;   // 4248 
           133 : coded = 13'b1000010111111;   // 4287 
           134 : coded = 13'b1000011000001;   // 4289 
           135 : coded = 13'b1000011100110;   // 4326 
           136 : coded = 13'b1000100000101;   // 4357 
           137 : coded = 13'b1000100100010;   // 4386 
           138 : coded = 13'b1000101011100;   // 4444 
           139 : coded = 13'b1000101111011;   // 4475 
           140 : coded = 13'b1000110001011;   // 4491 
           141 : coded = 13'b1000110101100;   // 4524 
           142 : coded = 13'b1000111010010;   // 4562 
           143 : coded = 13'b1000111110101;   // 4597 
           144 : coded = 13'b1001000001010;   // 4618 
           145 : coded = 13'b1001000101101;   // 4653 
           146 : coded = 13'b1001001010011;   // 4691 
           147 : coded = 13'b1001001110100;   // 4724 
           148 : coded = 13'b1001010000100;   // 4740 
           149 : coded = 13'b1001010100011;   // 4771 
           150 : coded = 13'b1001011011101;   // 4829 
           151 : coded = 13'b1001011111010;   // 4858 
           152 : coded = 13'b1001100011001;   // 4889 
           153 : coded = 13'b1001100111110;   // 4926 
           154 : coded = 13'b1001101000000;   // 4928 
           155 : coded = 13'b1001101100111;   // 4967 
           156 : coded = 13'b1001110010111;   // 5015 
           157 : coded = 13'b1001110110000;   // 5040 
           158 : coded = 13'b1001111001110;   // 5070 
           159 : coded = 13'b1001111101001;   // 5097 
           160 : coded = 13'b1010000011101;   // 5149 
           161 : coded = 13'b1010000111010;   // 5178 
           162 : coded = 13'b1010001000100;   // 5188 
           163 : coded = 13'b1010001100011;   // 5219 
           164 : coded = 13'b1010010010011;   // 5267 
           165 : coded = 13'b1010010110100;   // 5300 
           166 : coded = 13'b1010011001010;   // 5322 
           167 : coded = 13'b1010011101101;   // 5357 
           168 : coded = 13'b1010100001110;   // 5390 
           169 : coded = 13'b1010100101001;   // 5417 
           170 : coded = 13'b1010101010111;   // 5463 
           171 : coded = 13'b1010101110000;   // 5488 
           172 : coded = 13'b1010110000000;   // 5504 
           173 : coded = 13'b1010110100111;   // 5543 
           174 : coded = 13'b1010111011001;   // 5593 
           175 : coded = 13'b1010111111110;   // 5630 
           176 : coded = 13'b1011000000001;   // 5633 
           177 : coded = 13'b1011000100110;   // 5670 
           178 : coded = 13'b1011001011000;   // 5720 
           179 : coded = 13'b1011001111111;   // 5759 
           180 : coded = 13'b1011010001111;   // 5775 
           181 : coded = 13'b1011010101000;   // 5800 
           182 : coded = 13'b1011011010110;   // 5846 
           183 : coded = 13'b1011011110001;   // 5873 
           184 : coded = 13'b1011100010010;   // 5906 
           185 : coded = 13'b1011100110101;   // 5941 
           186 : coded = 13'b1011101001011;   // 5963 
           187 : coded = 13'b1011101101100;   // 5996 
           188 : coded = 13'b1011110011100;   // 6044 
           189 : coded = 13'b1011110111011;   // 6075 
           190 : coded = 13'b1011111000101;   // 6085 
           191 : coded = 13'b1011111100010;   // 6114 
           192 : coded = 13'b1100000000011;   // 6147 
           193 : coded = 13'b1100000100100;   // 6180 
           194 : coded = 13'b1100001011010;   // 6234 
           195 : coded = 13'b1100001111101;   // 6269 
           196 : coded = 13'b1100010001101;   // 6285 
           197 : coded = 13'b1100010101010;   // 6314 
           198 : coded = 13'b1100011010100;   // 6356 
           199 : coded = 13'b1100011110011;   // 6387 
           200 : coded = 13'b1100100010000;   // 6416 
           201 : coded = 13'b1100100110111;   // 6455 
           202 : coded = 13'b1100101001001;   // 6473 
           203 : coded = 13'b1100101101110;   // 6510 
           204 : coded = 13'b1100110011110;   // 6558 
           205 : coded = 13'b1100110111001;   // 6585 
           206 : coded = 13'b1100111000111;   // 6599 
           207 : coded = 13'b1100111100000;   // 6624 
           208 : coded = 13'b1101000011111;   // 6687 
           209 : coded = 13'b1101000111000;   // 6712 
           210 : coded = 13'b1101001000110;   // 6726 
           211 : coded = 13'b1101001100001;   // 6753 
           212 : coded = 13'b1101010010001;   // 6801 
           213 : coded = 13'b1101010110110;   // 6838 
           214 : coded = 13'b1101011001000;   // 6856 
           215 : coded = 13'b1101011101111;   // 6895 
           216 : coded = 13'b1101100001100;   // 6924 
           217 : coded = 13'b1101100101011;   // 6955 
           218 : coded = 13'b1101101010101;   // 6997 
           219 : coded = 13'b1101101110010;   // 7026 
           220 : coded = 13'b1101110000010;   // 7042 
           221 : coded = 13'b1101110100101;   // 7077 
           222 : coded = 13'b1101111011011;   // 7131 
           223 : coded = 13'b1101111111100;   // 7164 
           224 : coded = 13'b1110000001000;   // 7176 
           225 : coded = 13'b1110000101111;   // 7215 
           226 : coded = 13'b1110001010001;   // 7249 
           227 : coded = 13'b1110001110110;   // 7286 
           228 : coded = 13'b1110010000110;   // 7302 
           229 : coded = 13'b1110010100001;   // 7329 
           230 : coded = 13'b1110011011111;   // 7391 
           231 : coded = 13'b1110011111000;   // 7416 
           232 : coded = 13'b1110100011011;   // 7451 
           233 : coded = 13'b1110100111100;   // 7484 
           234 : coded = 13'b1110101000010;   // 7490 
           235 : coded = 13'b1110101100101;   // 7525 
           236 : coded = 13'b1110110010101;   // 7573 
           237 : coded = 13'b1110110110010;   // 7602 
           238 : coded = 13'b1110111001100;   // 7628 
           239 : coded = 13'b1110111101011;   // 7659 
           240 : coded = 13'b1111000010100;   // 7700 
           241 : coded = 13'b1111000110011;   // 7731 
           242 : coded = 13'b1111001001101;   // 7757 
           243 : coded = 13'b1111001101010;   // 7786 
           244 : coded = 13'b1111010011010;   // 7834 
           245 : coded = 13'b1111010111101;   // 7869 
           246 : coded = 13'b1111011000011;   // 7875 
           247 : coded = 13'b1111011100100;   // 7908 
           248 : coded = 13'b1111100000111;   // 7943 
           249 : coded = 13'b1111100100000;   // 7968 
           250 : coded = 13'b1111101011110;   // 8030 
           251 : coded = 13'b1111101111001;   // 8057 
           252 : coded = 13'b1111110001001;   // 8073 
           253 : coded = 13'b1111110101110;   // 8110 
           254 : coded = 13'b1111111010000;   // 8144 
           255 : coded = 13'b1111111110111;   // 8183 
           256 : coded = 13'b0000000000000;   // 0 
           257 : coded = 13'b0000000100111;   // 39 
           258 : coded = 13'b0000001011001;   // 89 
           259 : coded = 13'b0000001111110;   // 126 
           260 : coded = 13'b0000010001110;   // 142 
           261 : coded = 13'b0000010101001;   // 169 
           262 : coded = 13'b0000011010111;   // 215 
           263 : coded = 13'b0000011110000;   // 240 
           264 : coded = 13'b0000100010011;   // 275 
           265 : coded = 13'b0000100110100;   // 308 
           266 : coded = 13'b0000101001010;   // 330 
           267 : coded = 13'b0000101101101;   // 365 
           268 : coded = 13'b0000110011101;   // 413 
           269 : coded = 13'b0000110111010;   // 442 
           270 : coded = 13'b0000111000100;   // 452 
           271 : coded = 13'b0000111100011;   // 483 
           272 : coded = 13'b0001000011100;   // 540 
           273 : coded = 13'b0001000111011;   // 571 
           274 : coded = 13'b0001001000101;   // 581 
           275 : coded = 13'b0001001100010;   // 610 
           276 : coded = 13'b0001010010010;   // 658 
           277 : coded = 13'b0001010110101;   // 693 
           278 : coded = 13'b0001011001011;   // 715 
           279 : coded = 13'b0001011101100;   // 748 
           280 : coded = 13'b0001100001111;   // 783 
           281 : coded = 13'b0001100101000;   // 808 
           282 : coded = 13'b0001101010110;   // 854 
           283 : coded = 13'b0001101110001;   // 881 
           284 : coded = 13'b0001110000001;   // 897 
           285 : coded = 13'b0001110100110;   // 934 
           286 : coded = 13'b0001111011000;   // 984 
           287 : coded = 13'b0001111111111;   // 1023 
           288 : coded = 13'b0010000001011;   // 1035 
           289 : coded = 13'b0010000101100;   // 1068 
           290 : coded = 13'b0010001010010;   // 1106 
           291 : coded = 13'b0010001110101;   // 1141 
           292 : coded = 13'b0010010000101;   // 1157 
           293 : coded = 13'b0010010100010;   // 1186 
           294 : coded = 13'b0010011011100;   // 1244 
           295 : coded = 13'b0010011111011;   // 1275 
           296 : coded = 13'b0010100011000;   // 1304 
           297 : coded = 13'b0010100111111;   // 1343 
           298 : coded = 13'b0010101000001;   // 1345 
           299 : coded = 13'b0010101100110;   // 1382 
           300 : coded = 13'b0010110010110;   // 1430 
           301 : coded = 13'b0010110110001;   // 1457 
           302 : coded = 13'b0010111001111;   // 1487 
           303 : coded = 13'b0010111101000;   // 1512 
           304 : coded = 13'b0011000010111;   // 1559 
           305 : coded = 13'b0011000110000;   // 1584 
           306 : coded = 13'b0011001001110;   // 1614 
           307 : coded = 13'b0011001101001;   // 1641 
           308 : coded = 13'b0011010011001;   // 1689 
           309 : coded = 13'b0011010111110;   // 1726 
           310 : coded = 13'b0011011000000;   // 1728 
           311 : coded = 13'b0011011100111;   // 1767 
           312 : coded = 13'b0011100000100;   // 1796 
           313 : coded = 13'b0011100100011;   // 1827 
           314 : coded = 13'b0011101011101;   // 1885 
           315 : coded = 13'b0011101111010;   // 1914 
           316 : coded = 13'b0011110001010;   // 1930 
           317 : coded = 13'b0011110101101;   // 1965 
           318 : coded = 13'b0011111010011;   // 2003 
           319 : coded = 13'b0011111110100;   // 2036 
           320 : coded = 13'b0100000010101;   // 2069 
           321 : coded = 13'b0100000110010;   // 2098 
           322 : coded = 13'b0100001001100;   // 2124 
           323 : coded = 13'b0100001101011;   // 2155 
           324 : coded = 13'b0100010011011;   // 2203 
           325 : coded = 13'b0100010111100;   // 2236 
           326 : coded = 13'b0100011000010;   // 2242 
           327 : coded = 13'b0100011100101;   // 2277 
           328 : coded = 13'b0100100000110;   // 2310 
           329 : coded = 13'b0100100100001;   // 2337 
           330 : coded = 13'b0100101011111;   // 2399 
           331 : coded = 13'b0100101111000;   // 2424 
           332 : coded = 13'b0100110001000;   // 2440 
           333 : coded = 13'b0100110101111;   // 2479 
           334 : coded = 13'b0100111010001;   // 2513 
           335 : coded = 13'b0100111110110;   // 2550 
           336 : coded = 13'b0101000001001;   // 2569 
           337 : coded = 13'b0101000101110;   // 2606 
           338 : coded = 13'b0101001010000;   // 2640 
           339 : coded = 13'b0101001110111;   // 2679 
           340 : coded = 13'b0101010000111;   // 2695 
           341 : coded = 13'b0101010100000;   // 2720 
           342 : coded = 13'b0101011011110;   // 2782 
           343 : coded = 13'b0101011111001;   // 2809 
           344 : coded = 13'b0101100011010;   // 2842 
           345 : coded = 13'b0101100111101;   // 2877 
           346 : coded = 13'b0101101000011;   // 2883 
           347 : coded = 13'b0101101100100;   // 2916 
           348 : coded = 13'b0101110010100;   // 2964 
           349 : coded = 13'b0101110110011;   // 2995 
           350 : coded = 13'b0101111001101;   // 3021 
           351 : coded = 13'b0101111101010;   // 3050 
           352 : coded = 13'b0110000011110;   // 3102 
           353 : coded = 13'b0110000111001;   // 3129 
           354 : coded = 13'b0110001000111;   // 3143 
           355 : coded = 13'b0110001100000;   // 3168 
           356 : coded = 13'b0110010010000;   // 3216 
           357 : coded = 13'b0110010110111;   // 3255 
           358 : coded = 13'b0110011001001;   // 3273 
           359 : coded = 13'b0110011101110;   // 3310 
           360 : coded = 13'b0110100001101;   // 3341 
           361 : coded = 13'b0110100101010;   // 3370 
           362 : coded = 13'b0110101010100;   // 3412 
           363 : coded = 13'b0110101110011;   // 3443 
           364 : coded = 13'b0110110000011;   // 3459 
           365 : coded = 13'b0110110100100;   // 3492 
           366 : coded = 13'b0110111011010;   // 3546 
           367 : coded = 13'b0110111111101;   // 3581 
           368 : coded = 13'b0111000000010;   // 3586 
           369 : coded = 13'b0111000100101;   // 3621 
           370 : coded = 13'b0111001011011;   // 3675 
           371 : coded = 13'b0111001111100;   // 3708 
           372 : coded = 13'b0111010001100;   // 3724 
           373 : coded = 13'b0111010101011;   // 3755 
           374 : coded = 13'b0111011010101;   // 3797 
           375 : coded = 13'b0111011110010;   // 3826 
           376 : coded = 13'b0111100010001;   // 3857 
           377 : coded = 13'b0111100110110;   // 3894 
           378 : coded = 13'b0111101001000;   // 3912 
           379 : coded = 13'b0111101101111;   // 3951 
           380 : coded = 13'b0111110011111;   // 3999 
           381 : coded = 13'b0111110111000;   // 4024 
           382 : coded = 13'b0111111000110;   // 4038 
           383 : coded = 13'b0111111100001;   // 4065 
           384 : coded = 13'b1000000010110;   // 4118 
           385 : coded = 13'b1000000110001;   // 4145 
           386 : coded = 13'b1000001001111;   // 4175 
           387 : coded = 13'b1000001101000;   // 4200 
           388 : coded = 13'b1000010011000;   // 4248 
           389 : coded = 13'b1000010111111;   // 4287 
           390 : coded = 13'b1000011000001;   // 4289 
           391 : coded = 13'b1000011100110;   // 4326 
           392 : coded = 13'b1000100000101;   // 4357 
           393 : coded = 13'b1000100100010;   // 4386 
           394 : coded = 13'b1000101011100;   // 4444 
           395 : coded = 13'b1000101111011;   // 4475 
           396 : coded = 13'b1000110001011;   // 4491 
           397 : coded = 13'b1000110101100;   // 4524 
           398 : coded = 13'b1000111010010;   // 4562 
           399 : coded = 13'b1000111110101;   // 4597 
           400 : coded = 13'b1001000001010;   // 4618 
           401 : coded = 13'b1001000101101;   // 4653 
           402 : coded = 13'b1001001010011;   // 4691 
           403 : coded = 13'b1001001110100;   // 4724 
           404 : coded = 13'b1001010000100;   // 4740 
           405 : coded = 13'b1001010100011;   // 4771 
           406 : coded = 13'b1001011011101;   // 4829 
           407 : coded = 13'b1001011111010;   // 4858 
           408 : coded = 13'b1001100011001;   // 4889 
           409 : coded = 13'b1001100111110;   // 4926 
           410 : coded = 13'b1001101000000;   // 4928 
           411 : coded = 13'b1001101100111;   // 4967 
           412 : coded = 13'b1001110010111;   // 5015 
           413 : coded = 13'b1001110110000;   // 5040 
           414 : coded = 13'b1001111001110;   // 5070 
           415 : coded = 13'b1001111101001;   // 5097 
           416 : coded = 13'b1010000011101;   // 5149 
           417 : coded = 13'b1010000111010;   // 5178 
           418 : coded = 13'b1010001000100;   // 5188 
           419 : coded = 13'b1010001100011;   // 5219 
           420 : coded = 13'b1010010010011;   // 5267 
           421 : coded = 13'b1010010110100;   // 5300 
           422 : coded = 13'b1010011001010;   // 5322 
           423 : coded = 13'b1010011101101;   // 5357 
           424 : coded = 13'b1010100001110;   // 5390 
           425 : coded = 13'b1010100101001;   // 5417 
           426 : coded = 13'b1010101010111;   // 5463 
           427 : coded = 13'b1010101110000;   // 5488 
           428 : coded = 13'b1010110000000;   // 5504 
           429 : coded = 13'b1010110100111;   // 5543 
           430 : coded = 13'b1010111011001;   // 5593 
           431 : coded = 13'b1010111111110;   // 5630 
           432 : coded = 13'b1011000000001;   // 5633 
           433 : coded = 13'b1011000100110;   // 5670 
           434 : coded = 13'b1011001011000;   // 5720 
           435 : coded = 13'b1011001111111;   // 5759 
           436 : coded = 13'b1011010001111;   // 5775 
           437 : coded = 13'b1011010101000;   // 5800 
           438 : coded = 13'b1011011010110;   // 5846 
           439 : coded = 13'b1011011110001;   // 5873 
           440 : coded = 13'b1011100010010;   // 5906 
           441 : coded = 13'b1011100110101;   // 5941 
           442 : coded = 13'b1011101001011;   // 5963 
           443 : coded = 13'b1011101101100;   // 5996 
           444 : coded = 13'b1011110011100;   // 6044 
           445 : coded = 13'b1011110111011;   // 6075 
           446 : coded = 13'b1011111000101;   // 6085 
           447 : coded = 13'b1011111100010;   // 6114 
           448 : coded = 13'b1100000000011;   // 6147 
           449 : coded = 13'b1100000100100;   // 6180 
           450 : coded = 13'b1100001011010;   // 6234 
           451 : coded = 13'b1100001111101;   // 6269 
           452 : coded = 13'b1100010001101;   // 6285 
           453 : coded = 13'b1100010101010;   // 6314 
           454 : coded = 13'b1100011010100;   // 6356 
           455 : coded = 13'b1100011110011;   // 6387 
           456 : coded = 13'b1100100010000;   // 6416 
           457 : coded = 13'b1100100110111;   // 6455 
           458 : coded = 13'b1100101001001;   // 6473 
           459 : coded = 13'b1100101101110;   // 6510 
           460 : coded = 13'b1100110011110;   // 6558 
           461 : coded = 13'b1100110111001;   // 6585 
           462 : coded = 13'b1100111000111;   // 6599 
           463 : coded = 13'b1100111100000;   // 6624 
           464 : coded = 13'b1101000011111;   // 6687 
           465 : coded = 13'b1101000111000;   // 6712 
           466 : coded = 13'b1101001000110;   // 6726 
           467 : coded = 13'b1101001100001;   // 6753 
           468 : coded = 13'b1101010010001;   // 6801 
           469 : coded = 13'b1101010110110;   // 6838 
           470 : coded = 13'b1101011001000;   // 6856 
           471 : coded = 13'b1101011101111;   // 6895 
           472 : coded = 13'b1101100001100;   // 6924 
           473 : coded = 13'b1101100101011;   // 6955 
           474 : coded = 13'b1101101010101;   // 6997 
           475 : coded = 13'b1101101110010;   // 7026 
           476 : coded = 13'b1101110000010;   // 7042 
           477 : coded = 13'b1101110100101;   // 7077 
           478 : coded = 13'b1101111011011;   // 7131 
           479 : coded = 13'b1101111111100;   // 7164 
           480 : coded = 13'b1110000001000;   // 7176 
           481 : coded = 13'b1110000101111;   // 7215 
           482 : coded = 13'b1110001010001;   // 7249 
           483 : coded = 13'b1110001110110;   // 7286 
           484 : coded = 13'b1110010000110;   // 7302 
           485 : coded = 13'b1110010100001;   // 7329 
           486 : coded = 13'b1110011011111;   // 7391 
           487 : coded = 13'b1110011111000;   // 7416 
           488 : coded = 13'b1110100011011;   // 7451 
           489 : coded = 13'b1110100111100;   // 7484 
           490 : coded = 13'b1110101000010;   // 7490 
           491 : coded = 13'b1110101100101;   // 7525 
           492 : coded = 13'b1110110010101;   // 7573 
           493 : coded = 13'b1110110110010;   // 7602 
           494 : coded = 13'b1110111001100;   // 7628 
           495 : coded = 13'b1110111101011;   // 7659 
           496 : coded = 13'b1111000010100;   // 7700 
           497 : coded = 13'b1111000110011;   // 7731 
           498 : coded = 13'b1111001001101;   // 7757 
           499 : coded = 13'b1111001101010;   // 7786 
           500 : coded = 13'b1111010011010;   // 7834 
           501 : coded = 13'b1111010111101;   // 7869 
           502 : coded = 13'b1111011000011;   // 7875 
           503 : coded = 13'b1111011100100;   // 7908 
           504 : coded = 13'b1111100000111;   // 7943 
           505 : coded = 13'b1111100100000;   // 7968 
           506 : coded = 13'b1111101011110;   // 8030 
           507 : coded = 13'b1111101111001;   // 8057 
           508 : coded = 13'b1111110001001;   // 8073 
           509 : coded = 13'b1111110101110;   // 8110 
           510 : coded = 13'b1111111010000;   // 8144 
           511 : coded = 13'b1111111110111;   // 8183 
           512 : coded = 13'b0000000000000;   // 0 
           513 : coded = 13'b0000000100111;   // 39 
           514 : coded = 13'b0000001011001;   // 89 
           515 : coded = 13'b0000001111110;   // 126 
           516 : coded = 13'b0000010001110;   // 142 
           517 : coded = 13'b0000010101001;   // 169 
           518 : coded = 13'b0000011010111;   // 215 
           519 : coded = 13'b0000011110000;   // 240 
           520 : coded = 13'b0000100010011;   // 275 
           521 : coded = 13'b0000100110100;   // 308 
           522 : coded = 13'b0000101001010;   // 330 
           523 : coded = 13'b0000101101101;   // 365 
           524 : coded = 13'b0000110011101;   // 413 
           525 : coded = 13'b0000110111010;   // 442 
           526 : coded = 13'b0000111000100;   // 452 
           527 : coded = 13'b0000111100011;   // 483 
           528 : coded = 13'b0001000011100;   // 540 
           529 : coded = 13'b0001000111011;   // 571 
           530 : coded = 13'b0001001000101;   // 581 
           531 : coded = 13'b0001001100010;   // 610 
           532 : coded = 13'b0001010010010;   // 658 
           533 : coded = 13'b0001010110101;   // 693 
           534 : coded = 13'b0001011001011;   // 715 
           535 : coded = 13'b0001011101100;   // 748 
           536 : coded = 13'b0001100001111;   // 783 
           537 : coded = 13'b0001100101000;   // 808 
           538 : coded = 13'b0001101010110;   // 854 
           539 : coded = 13'b0001101110001;   // 881 
           540 : coded = 13'b0001110000001;   // 897 
           541 : coded = 13'b0001110100110;   // 934 
           542 : coded = 13'b0001111011000;   // 984 
           543 : coded = 13'b0001111111111;   // 1023 
           544 : coded = 13'b0010000001011;   // 1035 
           545 : coded = 13'b0010000101100;   // 1068 
           546 : coded = 13'b0010001010010;   // 1106 
           547 : coded = 13'b0010001110101;   // 1141 
           548 : coded = 13'b0010010000101;   // 1157 
           549 : coded = 13'b0010010100010;   // 1186 
           550 : coded = 13'b0010011011100;   // 1244 
           551 : coded = 13'b0010011111011;   // 1275 
           552 : coded = 13'b0010100011000;   // 1304 
           553 : coded = 13'b0010100111111;   // 1343 
           554 : coded = 13'b0010101000001;   // 1345 
           555 : coded = 13'b0010101100110;   // 1382 
           556 : coded = 13'b0010110010110;   // 1430 
           557 : coded = 13'b0010110110001;   // 1457 
           558 : coded = 13'b0010111001111;   // 1487 
           559 : coded = 13'b0010111101000;   // 1512 
           560 : coded = 13'b0011000010111;   // 1559 
           561 : coded = 13'b0011000110000;   // 1584 
           562 : coded = 13'b0011001001110;   // 1614 
           563 : coded = 13'b0011001101001;   // 1641 
           564 : coded = 13'b0011010011001;   // 1689 
           565 : coded = 13'b0011010111110;   // 1726 
           566 : coded = 13'b0011011000000;   // 1728 
           567 : coded = 13'b0011011100111;   // 1767 
           568 : coded = 13'b0011100000100;   // 1796 
           569 : coded = 13'b0011100100011;   // 1827 
           570 : coded = 13'b0011101011101;   // 1885 
           571 : coded = 13'b0011101111010;   // 1914 
           572 : coded = 13'b0011110001010;   // 1930 
           573 : coded = 13'b0011110101101;   // 1965 
           574 : coded = 13'b0011111010011;   // 2003 
           575 : coded = 13'b0011111110100;   // 2036 
           576 : coded = 13'b0100000010101;   // 2069 
           577 : coded = 13'b0100000110010;   // 2098 
           578 : coded = 13'b0100001001100;   // 2124 
           579 : coded = 13'b0100001101011;   // 2155 
           580 : coded = 13'b0100010011011;   // 2203 
           581 : coded = 13'b0100010111100;   // 2236 
           582 : coded = 13'b0100011000010;   // 2242 
           583 : coded = 13'b0100011100101;   // 2277 
           584 : coded = 13'b0100100000110;   // 2310 
           585 : coded = 13'b0100100100001;   // 2337 
           586 : coded = 13'b0100101011111;   // 2399 
           587 : coded = 13'b0100101111000;   // 2424 
           588 : coded = 13'b0100110001000;   // 2440 
           589 : coded = 13'b0100110101111;   // 2479 
           590 : coded = 13'b0100111010001;   // 2513 
           591 : coded = 13'b0100111110110;   // 2550 
           592 : coded = 13'b0101000001001;   // 2569 
           593 : coded = 13'b0101000101110;   // 2606 
           594 : coded = 13'b0101001010000;   // 2640 
           595 : coded = 13'b0101001110111;   // 2679 
           596 : coded = 13'b0101010000111;   // 2695 
           597 : coded = 13'b0101010100000;   // 2720 
           598 : coded = 13'b0101011011110;   // 2782 
           599 : coded = 13'b0101011111001;   // 2809 
           600 : coded = 13'b0101100011010;   // 2842 
           601 : coded = 13'b0101100111101;   // 2877 
           602 : coded = 13'b0101101000011;   // 2883 
           603 : coded = 13'b0101101100100;   // 2916 
           604 : coded = 13'b0101110010100;   // 2964 
           605 : coded = 13'b0101110110011;   // 2995 
           606 : coded = 13'b0101111001101;   // 3021 
           607 : coded = 13'b0101111101010;   // 3050 
           608 : coded = 13'b0110000011110;   // 3102 
           609 : coded = 13'b0110000111001;   // 3129 
           610 : coded = 13'b0110001000111;   // 3143 
           611 : coded = 13'b0110001100000;   // 3168 
           612 : coded = 13'b0110010010000;   // 3216 
           613 : coded = 13'b0110010110111;   // 3255 
           614 : coded = 13'b0110011001001;   // 3273 
           615 : coded = 13'b0110011101110;   // 3310 
           616 : coded = 13'b0110100001101;   // 3341 
           617 : coded = 13'b0110100101010;   // 3370 
           618 : coded = 13'b0110101010100;   // 3412 
           619 : coded = 13'b0110101110011;   // 3443 
           620 : coded = 13'b0110110000011;   // 3459 
           621 : coded = 13'b0110110100100;   // 3492 
           622 : coded = 13'b0110111011010;   // 3546 
           623 : coded = 13'b0110111111101;   // 3581 
           624 : coded = 13'b0111000000010;   // 3586 
           625 : coded = 13'b0111000100101;   // 3621 
           626 : coded = 13'b0111001011011;   // 3675 
           627 : coded = 13'b0111001111100;   // 3708 
           628 : coded = 13'b0111010001100;   // 3724 
           629 : coded = 13'b0111010101011;   // 3755 
           630 : coded = 13'b0111011010101;   // 3797 
           631 : coded = 13'b0111011110010;   // 3826 
           632 : coded = 13'b0111100010001;   // 3857 
           633 : coded = 13'b0111100110110;   // 3894 
           634 : coded = 13'b0111101001000;   // 3912 
           635 : coded = 13'b0111101101111;   // 3951 
           636 : coded = 13'b0111110011111;   // 3999 
           637 : coded = 13'b0111110111000;   // 4024 
           638 : coded = 13'b0111111000110;   // 4038 
           639 : coded = 13'b0111111100001;   // 4065 
           640 : coded = 13'b1000000010110;   // 4118 
           641 : coded = 13'b1000000110001;   // 4145 
           642 : coded = 13'b1000001001111;   // 4175 
           643 : coded = 13'b1000001101000;   // 4200 
           644 : coded = 13'b1000010011000;   // 4248 
           645 : coded = 13'b1000010111111;   // 4287 
           646 : coded = 13'b1000011000001;   // 4289 
           647 : coded = 13'b1000011100110;   // 4326 
           648 : coded = 13'b1000100000101;   // 4357 
           649 : coded = 13'b1000100100010;   // 4386 
           650 : coded = 13'b1000101011100;   // 4444 
           651 : coded = 13'b1000101111011;   // 4475 
           652 : coded = 13'b1000110001011;   // 4491 
           653 : coded = 13'b1000110101100;   // 4524 
           654 : coded = 13'b1000111010010;   // 4562 
           655 : coded = 13'b1000111110101;   // 4597 
           656 : coded = 13'b1001000001010;   // 4618 
           657 : coded = 13'b1001000101101;   // 4653 
           658 : coded = 13'b1001001010011;   // 4691 
           659 : coded = 13'b1001001110100;   // 4724 
           660 : coded = 13'b1001010000100;   // 4740 
           661 : coded = 13'b1001010100011;   // 4771 
           662 : coded = 13'b1001011011101;   // 4829 
           663 : coded = 13'b1001011111010;   // 4858 
           664 : coded = 13'b1001100011001;   // 4889 
           665 : coded = 13'b1001100111110;   // 4926 
           666 : coded = 13'b1001101000000;   // 4928 
           667 : coded = 13'b1001101100111;   // 4967 
           668 : coded = 13'b1001110010111;   // 5015 
           669 : coded = 13'b1001110110000;   // 5040 
           670 : coded = 13'b1001111001110;   // 5070 
           671 : coded = 13'b1001111101001;   // 5097 
           672 : coded = 13'b1010000011101;   // 5149 
           673 : coded = 13'b1010000111010;   // 5178 
           674 : coded = 13'b1010001000100;   // 5188 
           675 : coded = 13'b1010001100011;   // 5219 
           676 : coded = 13'b1010010010011;   // 5267 
           677 : coded = 13'b1010010110100;   // 5300 
           678 : coded = 13'b1010011001010;   // 5322 
           679 : coded = 13'b1010011101101;   // 5357 
           680 : coded = 13'b1010100001110;   // 5390 
           681 : coded = 13'b1010100101001;   // 5417 
           682 : coded = 13'b1010101010111;   // 5463 
           683 : coded = 13'b1010101110000;   // 5488 
           684 : coded = 13'b1010110000000;   // 5504 
           685 : coded = 13'b1010110100111;   // 5543 
           686 : coded = 13'b1010111011001;   // 5593 
           687 : coded = 13'b1010111111110;   // 5630 
           688 : coded = 13'b1011000000001;   // 5633 
           689 : coded = 13'b1011000100110;   // 5670 
           690 : coded = 13'b1011001011000;   // 5720 
           691 : coded = 13'b1011001111111;   // 5759 
           692 : coded = 13'b1011010001111;   // 5775 
           693 : coded = 13'b1011010101000;   // 5800 
           694 : coded = 13'b1011011010110;   // 5846 
           695 : coded = 13'b1011011110001;   // 5873 
           696 : coded = 13'b1011100010010;   // 5906 
           697 : coded = 13'b1011100110101;   // 5941 
           698 : coded = 13'b1011101001011;   // 5963 
           699 : coded = 13'b1011101101100;   // 5996 
           700 : coded = 13'b1011110011100;   // 6044 
           701 : coded = 13'b1011110111011;   // 6075 
           702 : coded = 13'b1011111000101;   // 6085 
           703 : coded = 13'b1011111100010;   // 6114 
           704 : coded = 13'b1100000000011;   // 6147 
           705 : coded = 13'b1100000100100;   // 6180 
           706 : coded = 13'b1100001011010;   // 6234 
           707 : coded = 13'b1100001111101;   // 6269 
           708 : coded = 13'b1100010001101;   // 6285 
           709 : coded = 13'b1100010101010;   // 6314 
           710 : coded = 13'b1100011010100;   // 6356 
           711 : coded = 13'b1100011110011;   // 6387 
           712 : coded = 13'b1100100010000;   // 6416 
           713 : coded = 13'b1100100110111;   // 6455 
           714 : coded = 13'b1100101001001;   // 6473 
           715 : coded = 13'b1100101101110;   // 6510 
           716 : coded = 13'b1100110011110;   // 6558 
           717 : coded = 13'b1100110111001;   // 6585 
           718 : coded = 13'b1100111000111;   // 6599 
           719 : coded = 13'b1100111100000;   // 6624 
           720 : coded = 13'b1101000011111;   // 6687 
           721 : coded = 13'b1101000111000;   // 6712 
           722 : coded = 13'b1101001000110;   // 6726 
           723 : coded = 13'b1101001100001;   // 6753 
           724 : coded = 13'b1101010010001;   // 6801 
           725 : coded = 13'b1101010110110;   // 6838 
           726 : coded = 13'b1101011001000;   // 6856 
           727 : coded = 13'b1101011101111;   // 6895 
           728 : coded = 13'b1101100001100;   // 6924 
           729 : coded = 13'b1101100101011;   // 6955 
           730 : coded = 13'b1101101010101;   // 6997 
           731 : coded = 13'b1101101110010;   // 7026 
           732 : coded = 13'b1101110000010;   // 7042 
           733 : coded = 13'b1101110100101;   // 7077 
           734 : coded = 13'b1101111011011;   // 7131 
           735 : coded = 13'b1101111111100;   // 7164 
           736 : coded = 13'b1110000001000;   // 7176 
           737 : coded = 13'b1110000101111;   // 7215 
           738 : coded = 13'b1110001010001;   // 7249 
           739 : coded = 13'b1110001110110;   // 7286 
           740 : coded = 13'b1110010000110;   // 7302 
           741 : coded = 13'b1110010100001;   // 7329 
           742 : coded = 13'b1110011011111;   // 7391 
           743 : coded = 13'b1110011111000;   // 7416 
           744 : coded = 13'b1110100011011;   // 7451 
           745 : coded = 13'b1110100111100;   // 7484 
           746 : coded = 13'b1110101000010;   // 7490 
           747 : coded = 13'b1110101100101;   // 7525 
           748 : coded = 13'b1110110010101;   // 7573 
           749 : coded = 13'b1110110110010;   // 7602 
           750 : coded = 13'b1110111001100;   // 7628 
           751 : coded = 13'b1110111101011;   // 7659 
           752 : coded = 13'b1111000010100;   // 7700 
           753 : coded = 13'b1111000110011;   // 7731 
           754 : coded = 13'b1111001001101;   // 7757 
           755 : coded = 13'b1111001101010;   // 7786 
           756 : coded = 13'b1111010011010;   // 7834 
           757 : coded = 13'b1111010111101;   // 7869 
           758 : coded = 13'b1111011000011;   // 7875 
           759 : coded = 13'b1111011100100;   // 7908 
           760 : coded = 13'b1111100000111;   // 7943 
           761 : coded = 13'b1111100100000;   // 7968 
           762 : coded = 13'b1111101011110;   // 8030 
           763 : coded = 13'b1111101111001;   // 8057 
           764 : coded = 13'b1111110001001;   // 8073 
           765 : coded = 13'b1111110101110;   // 8110 
           766 : coded = 13'b1111111010000;   // 8144 
           767 : coded = 13'b1111111110111;   // 8183 
           768 : coded = 13'b0000000000000;   // 0 
           769 : coded = 13'b0000000100111;   // 39 
           770 : coded = 13'b0000001011001;   // 89 
           771 : coded = 13'b0000001111110;   // 126 
           772 : coded = 13'b0000010001110;   // 142 
           773 : coded = 13'b0000010101001;   // 169 
           774 : coded = 13'b0000011010111;   // 215 
           775 : coded = 13'b0000011110000;   // 240 
           776 : coded = 13'b0000100010011;   // 275 
           777 : coded = 13'b0000100110100;   // 308 
           778 : coded = 13'b0000101001010;   // 330 
           779 : coded = 13'b0000101101101;   // 365 
           780 : coded = 13'b0000110011101;   // 413 
           781 : coded = 13'b0000110111010;   // 442 
           782 : coded = 13'b0000111000100;   // 452 
           783 : coded = 13'b0000111100011;   // 483 
           784 : coded = 13'b0001000011100;   // 540 
           785 : coded = 13'b0001000111011;   // 571 
           786 : coded = 13'b0001001000101;   // 581 
           787 : coded = 13'b0001001100010;   // 610 
           788 : coded = 13'b0001010010010;   // 658 
           789 : coded = 13'b0001010110101;   // 693 
           790 : coded = 13'b0001011001011;   // 715 
           791 : coded = 13'b0001011101100;   // 748 
           792 : coded = 13'b0001100001111;   // 783 
           793 : coded = 13'b0001100101000;   // 808 
           794 : coded = 13'b0001101010110;   // 854 
           795 : coded = 13'b0001101110001;   // 881 
           796 : coded = 13'b0001110000001;   // 897 
           797 : coded = 13'b0001110100110;   // 934 
           798 : coded = 13'b0001111011000;   // 984 
           799 : coded = 13'b0001111111111;   // 1023 
           800 : coded = 13'b0010000001011;   // 1035 
           801 : coded = 13'b0010000101100;   // 1068 
           802 : coded = 13'b0010001010010;   // 1106 
           803 : coded = 13'b0010001110101;   // 1141 
           804 : coded = 13'b0010010000101;   // 1157 
           805 : coded = 13'b0010010100010;   // 1186 
           806 : coded = 13'b0010011011100;   // 1244 
           807 : coded = 13'b0010011111011;   // 1275 
           808 : coded = 13'b0010100011000;   // 1304 
           809 : coded = 13'b0010100111111;   // 1343 
           810 : coded = 13'b0010101000001;   // 1345 
           811 : coded = 13'b0010101100110;   // 1382 
           812 : coded = 13'b0010110010110;   // 1430 
           813 : coded = 13'b0010110110001;   // 1457 
           814 : coded = 13'b0010111001111;   // 1487 
           815 : coded = 13'b0010111101000;   // 1512 
           816 : coded = 13'b0011000010111;   // 1559 
           817 : coded = 13'b0011000110000;   // 1584 
           818 : coded = 13'b0011001001110;   // 1614 
           819 : coded = 13'b0011001101001;   // 1641 
           820 : coded = 13'b0011010011001;   // 1689 
           821 : coded = 13'b0011010111110;   // 1726 
           822 : coded = 13'b0011011000000;   // 1728 
           823 : coded = 13'b0011011100111;   // 1767 
           824 : coded = 13'b0011100000100;   // 1796 
           825 : coded = 13'b0011100100011;   // 1827 
           826 : coded = 13'b0011101011101;   // 1885 
           827 : coded = 13'b0011101111010;   // 1914 
           828 : coded = 13'b0011110001010;   // 1930 
           829 : coded = 13'b0011110101101;   // 1965 
           830 : coded = 13'b0011111010011;   // 2003 
           831 : coded = 13'b0011111110100;   // 2036 
           832 : coded = 13'b0100000010101;   // 2069 
           833 : coded = 13'b0100000110010;   // 2098 
           834 : coded = 13'b0100001001100;   // 2124 
           835 : coded = 13'b0100001101011;   // 2155 
           836 : coded = 13'b0100010011011;   // 2203 
           837 : coded = 13'b0100010111100;   // 2236 
           838 : coded = 13'b0100011000010;   // 2242 
           839 : coded = 13'b0100011100101;   // 2277 
           840 : coded = 13'b0100100000110;   // 2310 
           841 : coded = 13'b0100100100001;   // 2337 
           842 : coded = 13'b0100101011111;   // 2399 
           843 : coded = 13'b0100101111000;   // 2424 
           844 : coded = 13'b0100110001000;   // 2440 
           845 : coded = 13'b0100110101111;   // 2479 
           846 : coded = 13'b0100111010001;   // 2513 
           847 : coded = 13'b0100111110110;   // 2550 
           848 : coded = 13'b0101000001001;   // 2569 
           849 : coded = 13'b0101000101110;   // 2606 
           850 : coded = 13'b0101001010000;   // 2640 
           851 : coded = 13'b0101001110111;   // 2679 
           852 : coded = 13'b0101010000111;   // 2695 
           853 : coded = 13'b0101010100000;   // 2720 
           854 : coded = 13'b0101011011110;   // 2782 
           855 : coded = 13'b0101011111001;   // 2809 
           856 : coded = 13'b0101100011010;   // 2842 
           857 : coded = 13'b0101100111101;   // 2877 
           858 : coded = 13'b0101101000011;   // 2883 
           859 : coded = 13'b0101101100100;   // 2916 
           860 : coded = 13'b0101110010100;   // 2964 
           861 : coded = 13'b0101110110011;   // 2995 
           862 : coded = 13'b0101111001101;   // 3021 
           863 : coded = 13'b0101111101010;   // 3050 
           864 : coded = 13'b0110000011110;   // 3102 
           865 : coded = 13'b0110000111001;   // 3129 
           866 : coded = 13'b0110001000111;   // 3143 
           867 : coded = 13'b0110001100000;   // 3168 
           868 : coded = 13'b0110010010000;   // 3216 
           869 : coded = 13'b0110010110111;   // 3255 
           870 : coded = 13'b0110011001001;   // 3273 
           871 : coded = 13'b0110011101110;   // 3310 
           872 : coded = 13'b0110100001101;   // 3341 
           873 : coded = 13'b0110100101010;   // 3370 
           874 : coded = 13'b0110101010100;   // 3412 
           875 : coded = 13'b0110101110011;   // 3443 
           876 : coded = 13'b0110110000011;   // 3459 
           877 : coded = 13'b0110110100100;   // 3492 
           878 : coded = 13'b0110111011010;   // 3546 
           879 : coded = 13'b0110111111101;   // 3581 
           880 : coded = 13'b0111000000010;   // 3586 
           881 : coded = 13'b0111000100101;   // 3621 
           882 : coded = 13'b0111001011011;   // 3675 
           883 : coded = 13'b0111001111100;   // 3708 
           884 : coded = 13'b0111010001100;   // 3724 
           885 : coded = 13'b0111010101011;   // 3755 
           886 : coded = 13'b0111011010101;   // 3797 
           887 : coded = 13'b0111011110010;   // 3826 
           888 : coded = 13'b0111100010001;   // 3857 
           889 : coded = 13'b0111100110110;   // 3894 
           890 : coded = 13'b0111101001000;   // 3912 
           891 : coded = 13'b0111101101111;   // 3951 
           892 : coded = 13'b0111110011111;   // 3999 
           893 : coded = 13'b0111110111000;   // 4024 
           894 : coded = 13'b0111111000110;   // 4038 
           895 : coded = 13'b0111111100001;   // 4065 
           896 : coded = 13'b1000000010110;   // 4118 
           897 : coded = 13'b1000000110001;   // 4145 
           898 : coded = 13'b1000001001111;   // 4175 
           899 : coded = 13'b1000001101000;   // 4200 
           900 : coded = 13'b1000010011000;   // 4248 
           901 : coded = 13'b1000010111111;   // 4287 
           902 : coded = 13'b1000011000001;   // 4289 
           903 : coded = 13'b1000011100110;   // 4326 
           904 : coded = 13'b1000100000101;   // 4357 
           905 : coded = 13'b1000100100010;   // 4386 
           906 : coded = 13'b1000101011100;   // 4444 
           907 : coded = 13'b1000101111011;   // 4475 
           908 : coded = 13'b1000110001011;   // 4491 
           909 : coded = 13'b1000110101100;   // 4524 
           910 : coded = 13'b1000111010010;   // 4562 
           911 : coded = 13'b1000111110101;   // 4597 
           912 : coded = 13'b1001000001010;   // 4618 
           913 : coded = 13'b1001000101101;   // 4653 
           914 : coded = 13'b1001001010011;   // 4691 
           915 : coded = 13'b1001001110100;   // 4724 
           916 : coded = 13'b1001010000100;   // 4740 
           917 : coded = 13'b1001010100011;   // 4771 
           918 : coded = 13'b1001011011101;   // 4829 
           919 : coded = 13'b1001011111010;   // 4858 
           920 : coded = 13'b1001100011001;   // 4889 
           921 : coded = 13'b1001100111110;   // 4926 
           922 : coded = 13'b1001101000000;   // 4928 
           923 : coded = 13'b1001101100111;   // 4967 
           924 : coded = 13'b1001110010111;   // 5015 
           925 : coded = 13'b1001110110000;   // 5040 
           926 : coded = 13'b1001111001110;   // 5070 
           927 : coded = 13'b1001111101001;   // 5097 
           928 : coded = 13'b1010000011101;   // 5149 
           929 : coded = 13'b1010000111010;   // 5178 
           930 : coded = 13'b1010001000100;   // 5188 
           931 : coded = 13'b1010001100011;   // 5219 
           932 : coded = 13'b1010010010011;   // 5267 
           933 : coded = 13'b1010010110100;   // 5300 
           934 : coded = 13'b1010011001010;   // 5322 
           935 : coded = 13'b1010011101101;   // 5357 
           936 : coded = 13'b1010100001110;   // 5390 
           937 : coded = 13'b1010100101001;   // 5417 
           938 : coded = 13'b1010101010111;   // 5463 
           939 : coded = 13'b1010101110000;   // 5488 
           940 : coded = 13'b1010110000000;   // 5504 
           941 : coded = 13'b1010110100111;   // 5543 
           942 : coded = 13'b1010111011001;   // 5593 
           943 : coded = 13'b1010111111110;   // 5630 
           944 : coded = 13'b1011000000001;   // 5633 
           945 : coded = 13'b1011000100110;   // 5670 
           946 : coded = 13'b1011001011000;   // 5720 
           947 : coded = 13'b1011001111111;   // 5759 
           948 : coded = 13'b1011010001111;   // 5775 
           949 : coded = 13'b1011010101000;   // 5800 
           950 : coded = 13'b1011011010110;   // 5846 
           951 : coded = 13'b1011011110001;   // 5873 
           952 : coded = 13'b1011100010010;   // 5906 
           953 : coded = 13'b1011100110101;   // 5941 
           954 : coded = 13'b1011101001011;   // 5963 
           955 : coded = 13'b1011101101100;   // 5996 
           956 : coded = 13'b1011110011100;   // 6044 
           957 : coded = 13'b1011110111011;   // 6075 
           958 : coded = 13'b1011111000101;   // 6085 
           959 : coded = 13'b1011111100010;   // 6114 
           960 : coded = 13'b1100000000011;   // 6147 
           961 : coded = 13'b1100000100100;   // 6180 
           962 : coded = 13'b1100001011010;   // 6234 
           963 : coded = 13'b1100001111101;   // 6269 
           964 : coded = 13'b1100010001101;   // 6285 
           965 : coded = 13'b1100010101010;   // 6314 
           966 : coded = 13'b1100011010100;   // 6356 
           967 : coded = 13'b1100011110011;   // 6387 
           968 : coded = 13'b1100100010000;   // 6416 
           969 : coded = 13'b1100100110111;   // 6455 
           970 : coded = 13'b1100101001001;   // 6473 
           971 : coded = 13'b1100101101110;   // 6510 
           972 : coded = 13'b1100110011110;   // 6558 
           973 : coded = 13'b1100110111001;   // 6585 
           974 : coded = 13'b1100111000111;   // 6599 
           975 : coded = 13'b1100111100000;   // 6624 
           976 : coded = 13'b1101000011111;   // 6687 
           977 : coded = 13'b1101000111000;   // 6712 
           978 : coded = 13'b1101001000110;   // 6726 
           979 : coded = 13'b1101001100001;   // 6753 
           980 : coded = 13'b1101010010001;   // 6801 
           981 : coded = 13'b1101010110110;   // 6838 
           982 : coded = 13'b1101011001000;   // 6856 
           983 : coded = 13'b1101011101111;   // 6895 
           984 : coded = 13'b1101100001100;   // 6924 
           985 : coded = 13'b1101100101011;   // 6955 
           986 : coded = 13'b1101101010101;   // 6997 
           987 : coded = 13'b1101101110010;   // 7026 
           988 : coded = 13'b1101110000010;   // 7042 
           989 : coded = 13'b1101110100101;   // 7077 
           990 : coded = 13'b1101111011011;   // 7131 
           991 : coded = 13'b1101111111100;   // 7164 
           992 : coded = 13'b1110000001000;   // 7176 
           993 : coded = 13'b1110000101111;   // 7215 
           994 : coded = 13'b1110001010001;   // 7249 
           995 : coded = 13'b1110001110110;   // 7286 
           996 : coded = 13'b1110010000110;   // 7302 
           997 : coded = 13'b1110010100001;   // 7329 
           998 : coded = 13'b1110011011111;   // 7391 
           999 : coded = 13'b1110011111000;   // 7416 
          1000 : coded = 13'b1110100011011;   // 7451 
          1001 : coded = 13'b1110100111100;   // 7484 
          1002 : coded = 13'b1110101000010;   // 7490 
          1003 : coded = 13'b1110101100101;   // 7525 
          1004 : coded = 13'b1110110010101;   // 7573 
          1005 : coded = 13'b1110110110010;   // 7602 
          1006 : coded = 13'b1110111001100;   // 7628 
          1007 : coded = 13'b1110111101011;   // 7659 
          1008 : coded = 13'b1111000010100;   // 7700 
          1009 : coded = 13'b1111000110011;   // 7731 
          1010 : coded = 13'b1111001001101;   // 7757 
          1011 : coded = 13'b1111001101010;   // 7786 
          1012 : coded = 13'b1111010011010;   // 7834 
          1013 : coded = 13'b1111010111101;   // 7869 
          1014 : coded = 13'b1111011000011;   // 7875 
          1015 : coded = 13'b1111011100100;   // 7908 
          1016 : coded = 13'b1111100000111;   // 7943 
          1017 : coded = 13'b1111100100000;   // 7968 
          1018 : coded = 13'b1111101011110;   // 8030 
          1019 : coded = 13'b1111101111001;   // 8057 
          1020 : coded = 13'b1111110001001;   // 8073 
          1021 : coded = 13'b1111110101110;   // 8110 
          1022 : coded = 13'b1111111010000;   // 8144 
          1023 : coded = 13'b1111111110111;   // 8183 
       default : coded = 13'bx; 
    endcase
endmodule
